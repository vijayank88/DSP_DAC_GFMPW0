// This is the unpowered netlist.
module DSP48 (user_clock2,
    wb_ACK,
    wb_CYC,
    wb_SEL,
    wb_STB,
    wb_WE,
    wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    wb_ADR,
    wb_DAT_MISO,
    wb_DAT_MOSI);
 input user_clock2;
 output wb_ACK;
 input wb_CYC;
 input wb_SEL;
 input wb_STB;
 input wb_WE;
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 input [31:0] wb_ADR;
 output [31:0] wb_DAT_MISO;
 input [31:0] wb_DAT_MOSI;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _zz_1_;
 wire \dacArea_dac_cnt_0[0] ;
 wire \dacArea_dac_cnt_0[1] ;
 wire \dacArea_dac_cnt_0[2] ;
 wire \dacArea_dac_cnt_0[3] ;
 wire \dacArea_dac_cnt_0[4] ;
 wire \dacArea_dac_cnt_0[5] ;
 wire \dacArea_dac_cnt_0[6] ;
 wire \dacArea_dac_cnt_1[0] ;
 wire \dacArea_dac_cnt_1[1] ;
 wire \dacArea_dac_cnt_1[2] ;
 wire \dacArea_dac_cnt_1[3] ;
 wire \dacArea_dac_cnt_1[4] ;
 wire \dacArea_dac_cnt_1[5] ;
 wire \dacArea_dac_cnt_1[6] ;
 wire \dacArea_dac_cnt_2[0] ;
 wire \dacArea_dac_cnt_2[1] ;
 wire \dacArea_dac_cnt_2[2] ;
 wire \dacArea_dac_cnt_2[3] ;
 wire \dacArea_dac_cnt_2[4] ;
 wire \dacArea_dac_cnt_2[5] ;
 wire \dacArea_dac_cnt_2[6] ;
 wire \dacArea_dac_cnt_3[0] ;
 wire \dacArea_dac_cnt_3[1] ;
 wire \dacArea_dac_cnt_3[2] ;
 wire \dacArea_dac_cnt_3[3] ;
 wire \dacArea_dac_cnt_3[4] ;
 wire \dacArea_dac_cnt_3[5] ;
 wire \dacArea_dac_cnt_3[6] ;
 wire \dacArea_dac_cnt_4[0] ;
 wire \dacArea_dac_cnt_4[1] ;
 wire \dacArea_dac_cnt_4[2] ;
 wire \dacArea_dac_cnt_4[3] ;
 wire \dacArea_dac_cnt_4[4] ;
 wire \dacArea_dac_cnt_4[5] ;
 wire \dacArea_dac_cnt_4[6] ;
 wire \dacArea_dac_cnt_5[0] ;
 wire \dacArea_dac_cnt_5[1] ;
 wire \dacArea_dac_cnt_5[2] ;
 wire \dacArea_dac_cnt_5[3] ;
 wire \dacArea_dac_cnt_5[4] ;
 wire \dacArea_dac_cnt_5[5] ;
 wire \dacArea_dac_cnt_5[6] ;
 wire \dacArea_dac_cnt_6[0] ;
 wire \dacArea_dac_cnt_6[1] ;
 wire \dacArea_dac_cnt_6[2] ;
 wire \dacArea_dac_cnt_6[3] ;
 wire \dacArea_dac_cnt_6[4] ;
 wire \dacArea_dac_cnt_6[5] ;
 wire \dacArea_dac_cnt_6[6] ;
 wire \dacArea_dac_cnt_7[0] ;
 wire \dacArea_dac_cnt_7[1] ;
 wire \dacArea_dac_cnt_7[2] ;
 wire \dacArea_dac_cnt_7[3] ;
 wire \dacArea_dac_cnt_7[4] ;
 wire \dacArea_dac_cnt_7[5] ;
 wire \dacArea_dac_cnt_7[6] ;
 wire \dspArea_regA[0] ;
 wire \dspArea_regA[10] ;
 wire \dspArea_regA[11] ;
 wire \dspArea_regA[12] ;
 wire \dspArea_regA[13] ;
 wire \dspArea_regA[14] ;
 wire \dspArea_regA[15] ;
 wire \dspArea_regA[16] ;
 wire \dspArea_regA[17] ;
 wire \dspArea_regA[18] ;
 wire \dspArea_regA[19] ;
 wire \dspArea_regA[1] ;
 wire \dspArea_regA[20] ;
 wire \dspArea_regA[21] ;
 wire \dspArea_regA[22] ;
 wire \dspArea_regA[23] ;
 wire \dspArea_regA[24] ;
 wire \dspArea_regA[2] ;
 wire \dspArea_regA[3] ;
 wire \dspArea_regA[4] ;
 wire \dspArea_regA[5] ;
 wire \dspArea_regA[6] ;
 wire \dspArea_regA[7] ;
 wire \dspArea_regA[8] ;
 wire \dspArea_regA[9] ;
 wire \dspArea_regB[0] ;
 wire \dspArea_regB[10] ;
 wire \dspArea_regB[11] ;
 wire \dspArea_regB[12] ;
 wire \dspArea_regB[13] ;
 wire \dspArea_regB[14] ;
 wire \dspArea_regB[15] ;
 wire \dspArea_regB[1] ;
 wire \dspArea_regB[2] ;
 wire \dspArea_regB[3] ;
 wire \dspArea_regB[4] ;
 wire \dspArea_regB[5] ;
 wire \dspArea_regB[6] ;
 wire \dspArea_regB[7] ;
 wire \dspArea_regB[8] ;
 wire \dspArea_regB[9] ;
 wire \dspArea_regP[0] ;
 wire \dspArea_regP[10] ;
 wire \dspArea_regP[11] ;
 wire \dspArea_regP[12] ;
 wire \dspArea_regP[13] ;
 wire \dspArea_regP[14] ;
 wire \dspArea_regP[15] ;
 wire \dspArea_regP[16] ;
 wire \dspArea_regP[17] ;
 wire \dspArea_regP[18] ;
 wire \dspArea_regP[19] ;
 wire \dspArea_regP[1] ;
 wire \dspArea_regP[20] ;
 wire \dspArea_regP[21] ;
 wire \dspArea_regP[22] ;
 wire \dspArea_regP[23] ;
 wire \dspArea_regP[24] ;
 wire \dspArea_regP[25] ;
 wire \dspArea_regP[26] ;
 wire \dspArea_regP[27] ;
 wire \dspArea_regP[28] ;
 wire \dspArea_regP[29] ;
 wire \dspArea_regP[2] ;
 wire \dspArea_regP[30] ;
 wire \dspArea_regP[31] ;
 wire \dspArea_regP[32] ;
 wire \dspArea_regP[33] ;
 wire \dspArea_regP[34] ;
 wire \dspArea_regP[35] ;
 wire \dspArea_regP[36] ;
 wire \dspArea_regP[37] ;
 wire \dspArea_regP[38] ;
 wire \dspArea_regP[39] ;
 wire \dspArea_regP[3] ;
 wire \dspArea_regP[40] ;
 wire \dspArea_regP[41] ;
 wire \dspArea_regP[42] ;
 wire \dspArea_regP[43] ;
 wire \dspArea_regP[44] ;
 wire \dspArea_regP[45] ;
 wire \dspArea_regP[46] ;
 wire \dspArea_regP[47] ;
 wire \dspArea_regP[4] ;
 wire \dspArea_regP[5] ;
 wire \dspArea_regP[6] ;
 wire \dspArea_regP[7] ;
 wire \dspArea_regP[8] ;
 wire \dspArea_regP[9] ;
 wire net231;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net232;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net233;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire clknet_0_wb_clk_i;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3709_ (.A1(net124),
    .A2(_zz_1_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3710_ (.I(_3265_),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3711_ (.A1(net83),
    .A2(net82),
    .A3(net85),
    .A4(net84),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3712_ (.A1(net79),
    .A2(net78),
    .A3(net81),
    .A4(net80),
    .Z(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3713_ (.A1(net74),
    .A2(net73),
    .A3(net76),
    .A4(net75),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3714_ (.A1(net87),
    .A2(net86),
    .A3(net90),
    .A4(net89),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _3715_ (.A1(_3267_),
    .A2(_3268_),
    .A3(_3269_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3716_ (.A1(_3266_),
    .A2(_3270_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3717_ (.A1(net70),
    .A2(net69),
    .A3(net72),
    .A4(net71),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3718_ (.A1(net97),
    .A2(net96),
    .A3(net68),
    .A4(net67),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3719_ (.A1(net77),
    .A2(net66),
    .A3(_3272_),
    .A4(_3273_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3720_ (.A1(_3271_),
    .A2(_3274_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3721_ (.I(net92),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3722_ (.A1(net93),
    .A2(net95),
    .A3(net94),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3723_ (.A1(_3276_),
    .A2(_3277_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3724_ (.A1(net88),
    .A2(_3278_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3725_ (.A1(net91),
    .A2(_3275_),
    .A3(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3726_ (.I(_3280_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3727_ (.I(net88),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3728_ (.I(net91),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3729_ (.A1(_3282_),
    .A2(_3283_),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3730_ (.A1(_3271_),
    .A2(_3274_),
    .A3(_3284_),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3731_ (.A1(net92),
    .A2(_3277_),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3732_ (.A1(_3285_),
    .A2(_3286_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3733_ (.I(_3287_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3734_ (.I(_3288_),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3735_ (.I(\dspArea_regA[0] ),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3736_ (.I(_3290_),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3737_ (.I(_3291_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3738_ (.I(_3292_),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3739_ (.I(_3293_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3740_ (.A1(_3282_),
    .A2(net91),
    .A3(_3275_),
    .A4(_3278_),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3741_ (.I(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3742_ (.I(_3296_),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3743_ (.A1(\dspArea_regP[32] ),
    .A2(_3281_),
    .B1(_3289_),
    .B2(_3294_),
    .C1(_3297_),
    .C2(\dspArea_regP[0] ),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3744_ (.I(_3298_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3745_ (.I(\dspArea_regA[1] ),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3746_ (.I(_3299_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3747_ (.I(_3300_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3748_ (.I(_3301_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3749_ (.A1(\dspArea_regP[33] ),
    .A2(_3281_),
    .B1(_3289_),
    .B2(_3302_),
    .C1(_3297_),
    .C2(\dspArea_regP[1] ),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3750_ (.I(_3303_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3751_ (.I(\dspArea_regA[2] ),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3752_ (.I(_3304_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3753_ (.I(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3754_ (.I(_3306_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3755_ (.I(_3307_),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3756_ (.A1(\dspArea_regP[34] ),
    .A2(_3281_),
    .B1(_3289_),
    .B2(_3308_),
    .C1(_3297_),
    .C2(\dspArea_regP[2] ),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3757_ (.I(_3309_),
    .ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3758_ (.I(_3287_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3759_ (.I(_3310_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3760_ (.I(\dspArea_regA[3] ),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3761_ (.I(_3312_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3762_ (.I(_3313_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3763_ (.I(_3314_),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3764_ (.I(_3315_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3765_ (.I(_3316_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_3296_),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3767_ (.A1(\dspArea_regP[35] ),
    .A2(_3281_),
    .B1(_3311_),
    .B2(_3317_),
    .C1(_3318_),
    .C2(\dspArea_regP[3] ),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3768_ (.I(_3319_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3769_ (.I(_3280_),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3770_ (.I(\dspArea_regA[4] ),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3771_ (.I(_3321_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3772_ (.I(_3322_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3773_ (.I(_3323_),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(_3324_),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3775_ (.I(_3325_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3776_ (.A1(\dspArea_regP[36] ),
    .A2(_3320_),
    .B1(_3311_),
    .B2(_3326_),
    .C1(_3318_),
    .C2(\dspArea_regP[4] ),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3777_ (.I(_3327_),
    .ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3778_ (.I(\dspArea_regA[5] ),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3779_ (.I(_3328_),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3780_ (.I(_3329_),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3781_ (.I(_3330_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3782_ (.I(_3331_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3783_ (.I(_3332_),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3784_ (.A1(\dspArea_regP[37] ),
    .A2(_3320_),
    .B1(_3311_),
    .B2(_3333_),
    .C1(_3318_),
    .C2(\dspArea_regP[5] ),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3785_ (.I(_3334_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3786_ (.I(\dspArea_regA[6] ),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3787_ (.I(_3335_),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3788_ (.I(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3789_ (.I(_3337_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3790_ (.I(_3338_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3791_ (.I(_3339_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3792_ (.A1(\dspArea_regP[38] ),
    .A2(_3320_),
    .B1(_3311_),
    .B2(_3340_),
    .C1(_3318_),
    .C2(\dspArea_regP[6] ),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3793_ (.I(_3341_),
    .ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3794_ (.I(_3288_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3795_ (.I(\dspArea_regA[7] ),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3796_ (.I(_3343_),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3797_ (.I(_3344_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3798_ (.I(_3345_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3799_ (.I(_3346_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3800_ (.I(_3347_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3801_ (.I(_3296_),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3802_ (.A1(\dspArea_regP[39] ),
    .A2(_3320_),
    .B1(_3342_),
    .B2(_3348_),
    .C1(_3349_),
    .C2(\dspArea_regP[7] ),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3803_ (.I(_3350_),
    .ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3804_ (.I(_3280_),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3805_ (.I(\dspArea_regA[8] ),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3806_ (.I(_3352_),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3807_ (.I(_3353_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3808_ (.I(_3354_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3809_ (.I(_3355_),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3810_ (.A1(\dspArea_regP[40] ),
    .A2(_3351_),
    .B1(_3342_),
    .B2(_3356_),
    .C1(_3349_),
    .C2(\dspArea_regP[8] ),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3811_ (.I(_3357_),
    .ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3812_ (.I(\dspArea_regA[9] ),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3813_ (.I(_3358_),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3814_ (.I(_3359_),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3815_ (.I(_3360_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3816_ (.I(_3361_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3817_ (.I(_3362_),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3818_ (.A1(\dspArea_regP[41] ),
    .A2(_3351_),
    .B1(_3342_),
    .B2(_3363_),
    .C1(_3349_),
    .C2(\dspArea_regP[9] ),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3819_ (.I(_3364_),
    .ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3820_ (.I(\dspArea_regP[42] ),
    .Z(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3821_ (.I(\dspArea_regA[10] ),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3822_ (.I(_3366_),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3823_ (.I(_3367_),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3824_ (.I(_3368_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3825_ (.I(_3369_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3826_ (.I(_3370_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3827_ (.A1(_3365_),
    .A2(_3351_),
    .B1(_3342_),
    .B2(_3371_),
    .C1(_3349_),
    .C2(\dspArea_regP[10] ),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3828_ (.I(_3372_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3829_ (.I(_3288_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3830_ (.I(\dspArea_regA[11] ),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3831_ (.I(_3374_),
    .Z(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3832_ (.I(_3375_),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3833_ (.I(_3376_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3834_ (.I(_3377_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3835_ (.I(_3378_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3836_ (.I(_3296_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3837_ (.A1(\dspArea_regP[43] ),
    .A2(_3351_),
    .B1(_3373_),
    .B2(_3379_),
    .C1(_3380_),
    .C2(\dspArea_regP[11] ),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3838_ (.I(_3381_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3839_ (.I(_3280_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3840_ (.I(\dspArea_regA[12] ),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3841_ (.I(_3383_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3842_ (.I(_3384_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3843_ (.I(_3385_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3844_ (.I(_3386_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3845_ (.A1(\dspArea_regP[44] ),
    .A2(_3382_),
    .B1(_3373_),
    .B2(_3387_),
    .C1(_3380_),
    .C2(\dspArea_regP[12] ),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3846_ (.I(_3388_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3847_ (.I(\dspArea_regA[13] ),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3848_ (.I(_3389_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3849_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3850_ (.I(_3391_),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3851_ (.I(_3392_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3852_ (.A1(\dspArea_regP[45] ),
    .A2(_3382_),
    .B1(_3373_),
    .B2(_3393_),
    .C1(_3380_),
    .C2(\dspArea_regP[13] ),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3853_ (.I(_3394_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3854_ (.I(\dspArea_regA[14] ),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3855_ (.I(_3395_),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3856_ (.I(_3396_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3857_ (.I(_3397_),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3858_ (.I(_3398_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3859_ (.I(_3399_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3860_ (.I(_3400_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3861_ (.A1(\dspArea_regP[46] ),
    .A2(_3382_),
    .B1(_3373_),
    .B2(_3401_),
    .C1(_3380_),
    .C2(\dspArea_regP[14] ),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3862_ (.I(_3402_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3863_ (.I(\dspArea_regA[15] ),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3864_ (.I(_3403_),
    .Z(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3865_ (.I(_3404_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3866_ (.I(_3405_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3867_ (.I(_3406_),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3868_ (.I(_3407_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3869_ (.I(_3408_),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3870_ (.I(_3409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3871_ (.I(_3295_),
    .Z(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3872_ (.A1(\dspArea_regP[47] ),
    .A2(_3382_),
    .B1(_3310_),
    .B2(_3410_),
    .C1(_3411_),
    .C2(\dspArea_regP[15] ),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3873_ (.I(_3412_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3874_ (.I(\dspArea_regA[16] ),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3875_ (.I(_3413_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3876_ (.I(_3414_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3877_ (.I(_3415_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3878_ (.I(_3416_),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3879_ (.I(_3310_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3880_ (.A1(_3417_),
    .A2(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3881_ (.I(_3411_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3882_ (.A1(\dspArea_regP[16] ),
    .A2(_3420_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3883_ (.A1(_3419_),
    .A2(_3421_),
    .ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3884_ (.I(\dspArea_regA[17] ),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3885_ (.I(_3422_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3886_ (.I(_3423_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3887_ (.I(_3424_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3888_ (.I(_3425_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3889_ (.I(_3426_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3890_ (.A1(_3427_),
    .A2(_3418_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3891_ (.I(_3411_),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3892_ (.A1(\dspArea_regP[17] ),
    .A2(_3429_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3893_ (.A1(_3428_),
    .A2(_3430_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3894_ (.I(\dspArea_regA[18] ),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3895_ (.I(_3431_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3896_ (.I(_3432_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3897_ (.I(_3433_),
    .Z(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3898_ (.I(_3434_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3899_ (.A1(_3435_),
    .A2(_3418_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3900_ (.A1(\dspArea_regP[18] ),
    .A2(_3429_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3901_ (.A1(_3436_),
    .A2(_3437_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3902_ (.I(\dspArea_regA[19] ),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3903_ (.I(_3438_),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3904_ (.I(_3439_),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3905_ (.I(_3440_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3906_ (.I(_3441_),
    .Z(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3907_ (.I(_3442_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3908_ (.I(_3443_),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3909_ (.A1(_3444_),
    .A2(_3418_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3910_ (.A1(\dspArea_regP[19] ),
    .A2(_3429_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3911_ (.A1(_3445_),
    .A2(_3446_),
    .ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3912_ (.I(\dspArea_regA[20] ),
    .Z(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3913_ (.I(_3447_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3914_ (.I(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3915_ (.I(_3449_),
    .Z(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3916_ (.I(_3450_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3917_ (.I(_3451_),
    .Z(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3918_ (.I(_3310_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3919_ (.A1(_3452_),
    .A2(_3453_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3920_ (.A1(\dspArea_regP[20] ),
    .A2(_3429_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3921_ (.A1(_3454_),
    .A2(_3455_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3922_ (.I(\dspArea_regA[21] ),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3923_ (.I(_3456_),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3924_ (.I(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3925_ (.I(_3458_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3926_ (.I(_3459_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3927_ (.I(_3460_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3928_ (.A1(_3461_),
    .A2(_3453_),
    .ZN(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3929_ (.I(_3411_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3930_ (.A1(\dspArea_regP[21] ),
    .A2(_3463_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3931_ (.A1(_3462_),
    .A2(_3464_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3932_ (.I(\dspArea_regA[22] ),
    .Z(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3933_ (.I(_3465_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3934_ (.I(_3466_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(_3467_),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3936_ (.I(_3468_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3937_ (.A1(_3469_),
    .A2(_3453_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3938_ (.A1(\dspArea_regP[22] ),
    .A2(_3463_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3939_ (.A1(_3470_),
    .A2(_3471_),
    .ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(\dspArea_regA[23] ),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3941_ (.I(_3472_),
    .Z(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3942_ (.I(_3473_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3943_ (.I(_3474_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3944_ (.A1(_3475_),
    .A2(_3453_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3945_ (.A1(\dspArea_regP[23] ),
    .A2(_3463_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3946_ (.A1(_3476_),
    .A2(_3477_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3947_ (.I(\dspArea_regA[24] ),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3948_ (.I(_3478_),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3949_ (.I(_3479_),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3950_ (.I(_3480_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3951_ (.I(_3481_),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3952_ (.I(_3482_),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3953_ (.A1(_3483_),
    .A2(_3289_),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3954_ (.A1(\dspArea_regP[24] ),
    .A2(_3463_),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3955_ (.A1(_3484_),
    .A2(_3485_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_3297_),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3957_ (.A1(\dspArea_regP[25] ),
    .A2(_3486_),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3958_ (.A1(\dspArea_regP[26] ),
    .A2(_3486_),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3959_ (.A1(\dspArea_regP[27] ),
    .A2(_3486_),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3960_ (.A1(\dspArea_regP[28] ),
    .A2(_3486_),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3961_ (.A1(\dspArea_regP[29] ),
    .A2(_3420_),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3962_ (.A1(\dspArea_regP[30] ),
    .A2(_3420_),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3963_ (.A1(\dspArea_regP[31] ),
    .A2(_3420_),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3964_ (.I(net126),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3965_ (.I(_3487_),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3966_ (.I(_3488_),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3967_ (.A1(net124),
    .A2(net98),
    .A3(_3489_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3968_ (.I(net126),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3969_ (.I(_3490_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3970_ (.I(_3491_),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3971_ (.A1(\dacArea_dac_cnt_0[0] ),
    .A2(net1),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3972_ (.A1(\dacArea_dac_cnt_0[0] ),
    .A2(net1),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3973_ (.A1(_3492_),
    .A2(_3493_),
    .A3(_3494_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3974_ (.A1(\dacArea_dac_cnt_0[1] ),
    .A2(net12),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3975_ (.A1(_3494_),
    .A2(_3495_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3976_ (.A1(_3494_),
    .A2(_3495_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3977_ (.A1(_3489_),
    .A2(_3496_),
    .A3(_3497_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3978_ (.I(_3488_),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3979_ (.I(_3498_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3980_ (.A1(\dacArea_dac_cnt_0[1] ),
    .A2(net12),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3981_ (.A1(_3500_),
    .A2(_3497_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3982_ (.A1(\dacArea_dac_cnt_0[2] ),
    .A2(net23),
    .A3(_3501_),
    .ZN(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3983_ (.A1(_3499_),
    .A2(_3502_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3984_ (.A1(\dacArea_dac_cnt_0[2] ),
    .A2(net23),
    .ZN(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3985_ (.A1(_3501_),
    .A2(_3503_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3986_ (.A1(\dacArea_dac_cnt_0[2] ),
    .A2(net23),
    .B(_3504_),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3987_ (.A1(\dacArea_dac_cnt_0[3] ),
    .A2(net34),
    .A3(_3505_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3988_ (.A1(_3499_),
    .A2(_3506_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3989_ (.A1(\dacArea_dac_cnt_0[3] ),
    .A2(net34),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3990_ (.A1(\dacArea_dac_cnt_0[3] ),
    .A2(net34),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3991_ (.A1(_3507_),
    .A2(_3505_),
    .B(_3508_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3992_ (.A1(\dacArea_dac_cnt_0[4] ),
    .A2(net45),
    .A3(_3509_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3993_ (.A1(_3499_),
    .A2(_3510_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3994_ (.A1(\dacArea_dac_cnt_0[4] ),
    .A2(net45),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3995_ (.A1(\dacArea_dac_cnt_0[4] ),
    .A2(net45),
    .B(_3509_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3996_ (.A1(_3511_),
    .A2(_3512_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3997_ (.A1(\dacArea_dac_cnt_0[5] ),
    .A2(net56),
    .A3(_3513_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3998_ (.A1(_3499_),
    .A2(_3514_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3999_ (.I(_3488_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4000_ (.I(_3515_),
    .Z(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4001_ (.A1(\dacArea_dac_cnt_0[5] ),
    .A2(net56),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4002_ (.A1(_3517_),
    .A2(_3513_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4003_ (.A1(\dacArea_dac_cnt_0[5] ),
    .A2(net56),
    .B(_3518_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4004_ (.A1(\dacArea_dac_cnt_0[6] ),
    .A2(net61),
    .A3(_3519_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4005_ (.A1(_3516_),
    .A2(_3520_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4006_ (.I(_3490_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4007_ (.I(_3521_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4008_ (.A1(\dacArea_dac_cnt_0[6] ),
    .A2(net61),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4009_ (.A1(\dacArea_dac_cnt_0[6] ),
    .A2(net61),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4010_ (.A1(_3523_),
    .A2(_3519_),
    .B(_3524_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4011_ (.A1(net199),
    .A2(net62),
    .A3(_3525_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4012_ (.A1(_3522_),
    .A2(_3526_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4013_ (.A1(\dacArea_dac_cnt_1[0] ),
    .A2(net63),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4014_ (.A1(\dacArea_dac_cnt_1[0] ),
    .A2(net63),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4015_ (.A1(_3492_),
    .A2(_3527_),
    .A3(_3528_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4016_ (.A1(\dacArea_dac_cnt_1[1] ),
    .A2(net64),
    .Z(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4017_ (.A1(_3528_),
    .A2(_3529_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4018_ (.A1(_3528_),
    .A2(_3529_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4019_ (.A1(_3489_),
    .A2(_3530_),
    .A3(_3531_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4020_ (.A1(\dacArea_dac_cnt_1[1] ),
    .A2(net64),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4021_ (.A1(_3532_),
    .A2(_3531_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4022_ (.A1(\dacArea_dac_cnt_1[2] ),
    .A2(net2),
    .A3(_3533_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4023_ (.A1(_3516_),
    .A2(_3534_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4024_ (.A1(\dacArea_dac_cnt_1[2] ),
    .A2(net2),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4025_ (.A1(_3533_),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4026_ (.A1(\dacArea_dac_cnt_1[2] ),
    .A2(net2),
    .B(_3536_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4027_ (.A1(\dacArea_dac_cnt_1[3] ),
    .A2(net3),
    .A3(_3537_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4028_ (.A1(_3516_),
    .A2(_3538_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4029_ (.A1(\dacArea_dac_cnt_1[3] ),
    .A2(net3),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4030_ (.A1(\dacArea_dac_cnt_1[3] ),
    .A2(net3),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4031_ (.A1(_3539_),
    .A2(_3537_),
    .B(_3540_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4032_ (.A1(\dacArea_dac_cnt_1[4] ),
    .A2(net4),
    .A3(_3541_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4033_ (.A1(_3516_),
    .A2(_3542_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4034_ (.I(_3515_),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4035_ (.A1(\dacArea_dac_cnt_1[4] ),
    .A2(net4),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4036_ (.A1(\dacArea_dac_cnt_1[4] ),
    .A2(net4),
    .B(_3541_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4037_ (.A1(_3544_),
    .A2(_3545_),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4038_ (.A1(\dacArea_dac_cnt_1[5] ),
    .A2(net5),
    .A3(_3546_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4039_ (.A1(_3543_),
    .A2(_3547_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4040_ (.A1(\dacArea_dac_cnt_1[5] ),
    .A2(net5),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4041_ (.A1(_3548_),
    .A2(_3546_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4042_ (.A1(\dacArea_dac_cnt_1[5] ),
    .A2(net5),
    .B(_3549_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4043_ (.A1(\dacArea_dac_cnt_1[6] ),
    .A2(net6),
    .A3(_3550_),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4044_ (.A1(_3543_),
    .A2(_3551_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4045_ (.A1(\dacArea_dac_cnt_1[6] ),
    .A2(net6),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4046_ (.A1(\dacArea_dac_cnt_1[6] ),
    .A2(net6),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4047_ (.A1(_3552_),
    .A2(_3550_),
    .B(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4048_ (.A1(net198),
    .A2(net7),
    .A3(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4049_ (.A1(_3522_),
    .A2(_3555_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4050_ (.A1(\dacArea_dac_cnt_2[0] ),
    .A2(net8),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4051_ (.A1(\dacArea_dac_cnt_2[0] ),
    .A2(net8),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4052_ (.A1(_3492_),
    .A2(_3556_),
    .A3(_3557_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4053_ (.I(_3487_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4054_ (.I(_3558_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4055_ (.A1(\dacArea_dac_cnt_2[1] ),
    .A2(net9),
    .Z(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4056_ (.A1(_3557_),
    .A2(_3560_),
    .Z(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4057_ (.A1(_3557_),
    .A2(_3560_),
    .ZN(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4058_ (.A1(_3559_),
    .A2(_3561_),
    .A3(_3562_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4059_ (.A1(\dacArea_dac_cnt_2[1] ),
    .A2(net9),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4060_ (.A1(_3563_),
    .A2(_3562_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4061_ (.A1(\dacArea_dac_cnt_2[2] ),
    .A2(net10),
    .A3(_3564_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4062_ (.A1(_3543_),
    .A2(_3565_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4063_ (.A1(\dacArea_dac_cnt_2[2] ),
    .A2(net10),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4064_ (.A1(_3564_),
    .A2(_3566_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4065_ (.A1(\dacArea_dac_cnt_2[2] ),
    .A2(net10),
    .B(_3567_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4066_ (.A1(\dacArea_dac_cnt_2[3] ),
    .A2(net11),
    .A3(_3568_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4067_ (.A1(_3543_),
    .A2(_3569_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4068_ (.I(_3515_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4069_ (.A1(\dacArea_dac_cnt_2[3] ),
    .A2(net11),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4070_ (.A1(\dacArea_dac_cnt_2[3] ),
    .A2(net11),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4071_ (.A1(_3571_),
    .A2(_3568_),
    .B(_3572_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4072_ (.A1(\dacArea_dac_cnt_2[4] ),
    .A2(net13),
    .A3(_3573_),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4073_ (.A1(_3570_),
    .A2(_3574_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4074_ (.A1(\dacArea_dac_cnt_2[4] ),
    .A2(net13),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4075_ (.A1(\dacArea_dac_cnt_2[4] ),
    .A2(net13),
    .B(_3573_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4076_ (.A1(_3575_),
    .A2(_3576_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4077_ (.A1(\dacArea_dac_cnt_2[5] ),
    .A2(net14),
    .A3(_3577_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4078_ (.A1(_3570_),
    .A2(_3578_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4079_ (.A1(\dacArea_dac_cnt_2[5] ),
    .A2(net14),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4080_ (.A1(_3579_),
    .A2(_3577_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4081_ (.A1(\dacArea_dac_cnt_2[5] ),
    .A2(net14),
    .B(_3580_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4082_ (.A1(\dacArea_dac_cnt_2[6] ),
    .A2(net15),
    .A3(_3581_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4083_ (.A1(_3570_),
    .A2(_3582_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4084_ (.A1(\dacArea_dac_cnt_2[6] ),
    .A2(net15),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4085_ (.A1(\dacArea_dac_cnt_2[6] ),
    .A2(net15),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4086_ (.A1(_3583_),
    .A2(_3581_),
    .B(_3584_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4087_ (.A1(net197),
    .A2(net16),
    .A3(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4088_ (.A1(_3522_),
    .A2(_3586_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4089_ (.I(_3491_),
    .Z(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4090_ (.A1(\dacArea_dac_cnt_3[0] ),
    .A2(net17),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4091_ (.A1(\dacArea_dac_cnt_3[0] ),
    .A2(net17),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4092_ (.A1(_3587_),
    .A2(_3588_),
    .A3(_3589_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4093_ (.A1(\dacArea_dac_cnt_3[1] ),
    .A2(net18),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4094_ (.A1(_3589_),
    .A2(_3590_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4095_ (.A1(_3589_),
    .A2(_3590_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4096_ (.A1(_3559_),
    .A2(_3591_),
    .A3(_3592_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4097_ (.A1(\dacArea_dac_cnt_3[1] ),
    .A2(net18),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4098_ (.A1(_3593_),
    .A2(_3592_),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4099_ (.A1(\dacArea_dac_cnt_3[2] ),
    .A2(net19),
    .A3(_3594_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4100_ (.A1(_3570_),
    .A2(_3595_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4101_ (.I(_3515_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4102_ (.A1(\dacArea_dac_cnt_3[2] ),
    .A2(net19),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4103_ (.A1(_3594_),
    .A2(_3597_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4104_ (.A1(\dacArea_dac_cnt_3[2] ),
    .A2(net19),
    .B(_3598_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4105_ (.A1(\dacArea_dac_cnt_3[3] ),
    .A2(net20),
    .A3(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4106_ (.A1(_3596_),
    .A2(_3600_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4107_ (.A1(\dacArea_dac_cnt_3[3] ),
    .A2(net20),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4108_ (.A1(\dacArea_dac_cnt_3[3] ),
    .A2(net20),
    .ZN(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4109_ (.A1(_3601_),
    .A2(_3599_),
    .B(_3602_),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4110_ (.A1(\dacArea_dac_cnt_3[4] ),
    .A2(net21),
    .A3(_3603_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4111_ (.A1(_3596_),
    .A2(_3604_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4112_ (.A1(\dacArea_dac_cnt_3[4] ),
    .A2(net21),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4113_ (.A1(\dacArea_dac_cnt_3[4] ),
    .A2(net21),
    .B(_3603_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4114_ (.A1(_3605_),
    .A2(_3606_),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4115_ (.A1(\dacArea_dac_cnt_3[5] ),
    .A2(net22),
    .A3(_3607_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4116_ (.A1(_3596_),
    .A2(_3608_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4117_ (.A1(\dacArea_dac_cnt_3[5] ),
    .A2(net22),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4118_ (.A1(_3609_),
    .A2(_3607_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4119_ (.A1(\dacArea_dac_cnt_3[5] ),
    .A2(net22),
    .B(_3610_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4120_ (.A1(\dacArea_dac_cnt_3[6] ),
    .A2(net24),
    .A3(_3611_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4121_ (.A1(_3596_),
    .A2(_3612_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4122_ (.A1(\dacArea_dac_cnt_3[6] ),
    .A2(net24),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4123_ (.A1(\dacArea_dac_cnt_3[6] ),
    .A2(net24),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4124_ (.A1(_3613_),
    .A2(_3611_),
    .B(_3614_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4125_ (.A1(net196),
    .A2(net25),
    .A3(_3615_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4126_ (.A1(_3522_),
    .A2(_3616_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4127_ (.A1(\dacArea_dac_cnt_4[0] ),
    .A2(net26),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4128_ (.A1(\dacArea_dac_cnt_4[0] ),
    .A2(net26),
    .Z(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4129_ (.A1(_3587_),
    .A2(_3617_),
    .A3(_3618_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4130_ (.A1(\dacArea_dac_cnt_4[1] ),
    .A2(net27),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4131_ (.A1(_3618_),
    .A2(_3619_),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4132_ (.A1(_3618_),
    .A2(_3619_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4133_ (.A1(_3559_),
    .A2(_3620_),
    .A3(_3621_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4134_ (.I(_3488_),
    .Z(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4135_ (.I(_3622_),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4136_ (.A1(\dacArea_dac_cnt_4[1] ),
    .A2(net27),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4137_ (.A1(_3624_),
    .A2(_3621_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4138_ (.A1(\dacArea_dac_cnt_4[2] ),
    .A2(net28),
    .A3(_3625_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4139_ (.A1(_3623_),
    .A2(_3626_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4140_ (.A1(\dacArea_dac_cnt_4[2] ),
    .A2(net28),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4141_ (.A1(_3625_),
    .A2(_3627_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4142_ (.A1(\dacArea_dac_cnt_4[2] ),
    .A2(net28),
    .B(_3628_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4143_ (.A1(\dacArea_dac_cnt_4[3] ),
    .A2(net29),
    .A3(_3629_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4144_ (.A1(_3623_),
    .A2(_3630_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4145_ (.A1(\dacArea_dac_cnt_4[3] ),
    .A2(net29),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4146_ (.A1(\dacArea_dac_cnt_4[3] ),
    .A2(net29),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4147_ (.A1(_3631_),
    .A2(_3629_),
    .B(_3632_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4148_ (.A1(\dacArea_dac_cnt_4[4] ),
    .A2(net30),
    .A3(_3633_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4149_ (.A1(_3623_),
    .A2(_3634_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4150_ (.A1(\dacArea_dac_cnt_4[4] ),
    .A2(net30),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4151_ (.A1(\dacArea_dac_cnt_4[4] ),
    .A2(net30),
    .B(_3633_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4152_ (.A1(_3635_),
    .A2(_3636_),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4153_ (.A1(\dacArea_dac_cnt_4[5] ),
    .A2(net31),
    .A3(_3637_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4154_ (.A1(_3623_),
    .A2(_3638_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4155_ (.I(_3622_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4156_ (.A1(\dacArea_dac_cnt_4[5] ),
    .A2(net31),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4157_ (.A1(\dacArea_dac_cnt_4[5] ),
    .A2(net31),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4158_ (.A1(_3640_),
    .A2(_3637_),
    .B(_3641_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4159_ (.I(_3642_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4160_ (.A1(\dacArea_dac_cnt_4[6] ),
    .A2(net32),
    .A3(_3643_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4161_ (.A1(_3639_),
    .A2(_3644_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4162_ (.I(_3491_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4163_ (.A1(\dacArea_dac_cnt_4[6] ),
    .A2(net32),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4164_ (.A1(\dacArea_dac_cnt_4[6] ),
    .A2(net32),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4165_ (.A1(_3646_),
    .A2(_3643_),
    .B(_3647_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4166_ (.A1(net195),
    .A2(net33),
    .A3(_3648_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4167_ (.A1(_3645_),
    .A2(_3649_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4168_ (.A1(\dacArea_dac_cnt_5[0] ),
    .A2(net35),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4169_ (.A1(\dacArea_dac_cnt_5[0] ),
    .A2(net35),
    .Z(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4170_ (.A1(_3587_),
    .A2(_3650_),
    .A3(_3651_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4171_ (.A1(\dacArea_dac_cnt_5[1] ),
    .A2(net36),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4172_ (.A1(_3651_),
    .A2(_3652_),
    .Z(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4173_ (.A1(_3651_),
    .A2(_3652_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4174_ (.A1(_3559_),
    .A2(_3653_),
    .A3(_3654_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4175_ (.A1(\dacArea_dac_cnt_5[1] ),
    .A2(net36),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4176_ (.A1(_3655_),
    .A2(_3654_),
    .Z(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4177_ (.A1(\dacArea_dac_cnt_5[2] ),
    .A2(net37),
    .A3(_3656_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4178_ (.A1(_3639_),
    .A2(_3657_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4179_ (.A1(\dacArea_dac_cnt_5[2] ),
    .A2(net37),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4180_ (.A1(_3656_),
    .A2(_3658_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4181_ (.A1(\dacArea_dac_cnt_5[2] ),
    .A2(net37),
    .B(_3659_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4182_ (.A1(\dacArea_dac_cnt_5[3] ),
    .A2(net38),
    .A3(_3660_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4183_ (.A1(_3639_),
    .A2(_3661_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4184_ (.A1(\dacArea_dac_cnt_5[3] ),
    .A2(net38),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4185_ (.A1(\dacArea_dac_cnt_5[3] ),
    .A2(net38),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4186_ (.A1(_3662_),
    .A2(_3660_),
    .B(_3663_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4187_ (.A1(\dacArea_dac_cnt_5[4] ),
    .A2(net39),
    .A3(_3664_),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4188_ (.A1(_3639_),
    .A2(_3665_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4189_ (.I(_3622_),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4190_ (.A1(\dacArea_dac_cnt_5[4] ),
    .A2(net39),
    .ZN(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4191_ (.A1(\dacArea_dac_cnt_5[4] ),
    .A2(net39),
    .B(_3664_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4192_ (.A1(_3667_),
    .A2(_3668_),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4193_ (.A1(\dacArea_dac_cnt_5[5] ),
    .A2(net40),
    .A3(_3669_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4194_ (.A1(_3666_),
    .A2(_3670_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4195_ (.A1(\dacArea_dac_cnt_5[5] ),
    .A2(net40),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4196_ (.A1(_3671_),
    .A2(_3669_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4197_ (.A1(\dacArea_dac_cnt_5[5] ),
    .A2(net40),
    .B(_3672_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4198_ (.A1(\dacArea_dac_cnt_5[6] ),
    .A2(net41),
    .A3(_3673_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4199_ (.A1(_3666_),
    .A2(_3674_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4200_ (.A1(\dacArea_dac_cnt_5[6] ),
    .A2(net41),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4201_ (.A1(\dacArea_dac_cnt_5[6] ),
    .A2(net41),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4202_ (.A1(_3675_),
    .A2(_3673_),
    .B(_3676_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4203_ (.A1(net194),
    .A2(net42),
    .A3(_3677_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4204_ (.A1(_3645_),
    .A2(_3678_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4205_ (.A1(\dacArea_dac_cnt_6[0] ),
    .A2(net43),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4206_ (.A1(\dacArea_dac_cnt_6[0] ),
    .A2(net43),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4207_ (.A1(_3587_),
    .A2(_3679_),
    .A3(_3680_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4208_ (.I(_3558_),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4209_ (.A1(\dacArea_dac_cnt_6[1] ),
    .A2(net44),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4210_ (.A1(_3680_),
    .A2(_3682_),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4211_ (.A1(_3680_),
    .A2(_3682_),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4212_ (.A1(_3681_),
    .A2(_3683_),
    .A3(_3684_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4213_ (.A1(\dacArea_dac_cnt_6[1] ),
    .A2(net44),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4214_ (.A1(_3685_),
    .A2(_3684_),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4215_ (.A1(\dacArea_dac_cnt_6[2] ),
    .A2(net46),
    .A3(_3686_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4216_ (.A1(_3666_),
    .A2(_3687_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4217_ (.A1(\dacArea_dac_cnt_6[2] ),
    .A2(net46),
    .ZN(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4218_ (.A1(_3686_),
    .A2(_3688_),
    .ZN(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4219_ (.A1(\dacArea_dac_cnt_6[2] ),
    .A2(net46),
    .B(_3689_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4220_ (.A1(\dacArea_dac_cnt_6[3] ),
    .A2(net47),
    .A3(_3690_),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4221_ (.A1(_3666_),
    .A2(_3691_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4222_ (.I(_3622_),
    .Z(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4223_ (.A1(\dacArea_dac_cnt_6[3] ),
    .A2(net47),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4224_ (.A1(\dacArea_dac_cnt_6[3] ),
    .A2(net47),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4225_ (.A1(_3693_),
    .A2(_3690_),
    .B(_3694_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4226_ (.A1(\dacArea_dac_cnt_6[4] ),
    .A2(net48),
    .A3(_3695_),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4227_ (.A1(_3692_),
    .A2(_3696_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4228_ (.A1(\dacArea_dac_cnt_6[4] ),
    .A2(net48),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4229_ (.A1(\dacArea_dac_cnt_6[4] ),
    .A2(net48),
    .B(_3695_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4230_ (.A1(_3697_),
    .A2(_3698_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4231_ (.A1(\dacArea_dac_cnt_6[5] ),
    .A2(net49),
    .A3(_3699_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4232_ (.A1(_3692_),
    .A2(_3700_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4233_ (.A1(\dacArea_dac_cnt_6[5] ),
    .A2(net49),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4234_ (.A1(_3701_),
    .A2(_3699_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4235_ (.A1(\dacArea_dac_cnt_6[5] ),
    .A2(net49),
    .B(_3702_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4236_ (.A1(\dacArea_dac_cnt_6[6] ),
    .A2(net50),
    .A3(_3703_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4237_ (.A1(_3692_),
    .A2(_3704_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4238_ (.A1(\dacArea_dac_cnt_6[6] ),
    .A2(net50),
    .ZN(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4239_ (.A1(\dacArea_dac_cnt_6[6] ),
    .A2(net50),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4240_ (.A1(_3705_),
    .A2(_3703_),
    .B(_3706_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4241_ (.A1(net193),
    .A2(net51),
    .A3(_3707_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4242_ (.A1(_3645_),
    .A2(_3708_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4243_ (.I(_3491_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4244_ (.A1(\dacArea_dac_cnt_7[0] ),
    .A2(net52),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4245_ (.A1(\dacArea_dac_cnt_7[0] ),
    .A2(net52),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4246_ (.A1(_0154_),
    .A2(_0155_),
    .A3(_0156_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4247_ (.A1(\dacArea_dac_cnt_7[1] ),
    .A2(net53),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4248_ (.A1(_0156_),
    .A2(_0157_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4249_ (.A1(_0156_),
    .A2(_0157_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4250_ (.A1(_3681_),
    .A2(_0158_),
    .A3(_0159_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4251_ (.A1(\dacArea_dac_cnt_7[1] ),
    .A2(net53),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4252_ (.A1(_0160_),
    .A2(_0159_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4253_ (.A1(\dacArea_dac_cnt_7[2] ),
    .A2(net54),
    .A3(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4254_ (.A1(_3692_),
    .A2(_0162_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4255_ (.I(_3487_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4256_ (.I(_0163_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4257_ (.A1(\dacArea_dac_cnt_7[2] ),
    .A2(net54),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4258_ (.A1(_0161_),
    .A2(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4259_ (.A1(\dacArea_dac_cnt_7[2] ),
    .A2(net54),
    .B(_0166_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4260_ (.A1(\dacArea_dac_cnt_7[3] ),
    .A2(net55),
    .A3(_0167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4261_ (.A1(_0164_),
    .A2(_0168_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4262_ (.A1(\dacArea_dac_cnt_7[3] ),
    .A2(net55),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4263_ (.A1(\dacArea_dac_cnt_7[3] ),
    .A2(net55),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4264_ (.A1(_0169_),
    .A2(_0167_),
    .B(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4265_ (.A1(\dacArea_dac_cnt_7[4] ),
    .A2(net57),
    .A3(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4266_ (.A1(_0164_),
    .A2(_0172_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4267_ (.A1(\dacArea_dac_cnt_7[4] ),
    .A2(net57),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4268_ (.A1(\dacArea_dac_cnt_7[4] ),
    .A2(net57),
    .B(_0171_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4269_ (.A1(_0173_),
    .A2(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4270_ (.A1(\dacArea_dac_cnt_7[5] ),
    .A2(net58),
    .A3(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4271_ (.A1(_0164_),
    .A2(_0176_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4272_ (.A1(\dacArea_dac_cnt_7[5] ),
    .A2(net58),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4273_ (.A1(_0177_),
    .A2(_0175_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4274_ (.A1(\dacArea_dac_cnt_7[5] ),
    .A2(net58),
    .B(_0178_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4275_ (.A1(\dacArea_dac_cnt_7[6] ),
    .A2(net59),
    .A3(_0179_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4276_ (.A1(_0164_),
    .A2(_0180_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4277_ (.A1(\dacArea_dac_cnt_7[6] ),
    .A2(net59),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4278_ (.A1(\dacArea_dac_cnt_7[6] ),
    .A2(net59),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4279_ (.A1(_0181_),
    .A2(_0179_),
    .B(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4280_ (.A1(net192),
    .A2(net60),
    .A3(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4281_ (.A1(_3645_),
    .A2(_0184_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4282_ (.I(net99),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4283_ (.A1(net98),
    .A2(net125),
    .A3(net159),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4284_ (.A1(_3278_),
    .A2(_3285_),
    .A3(_0186_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4285_ (.I(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4286_ (.I(_0188_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4287_ (.I(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4288_ (.I(_0188_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4289_ (.A1(_3294_),
    .A2(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4290_ (.I(net126),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4291_ (.I(_0193_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4292_ (.A1(_0185_),
    .A2(_0190_),
    .B(_0192_),
    .C(_0194_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4293_ (.I(net110),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4294_ (.A1(_3302_),
    .A2(_0191_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4295_ (.A1(_0195_),
    .A2(_0190_),
    .B(_0196_),
    .C(_0194_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4296_ (.I(net116),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4297_ (.A1(_3308_),
    .A2(_0191_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4298_ (.A1(_0197_),
    .A2(_0190_),
    .B(_0198_),
    .C(_0194_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4299_ (.I(net117),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4300_ (.I(_0187_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4301_ (.I(_0200_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4302_ (.A1(_3317_),
    .A2(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4303_ (.A1(_0199_),
    .A2(_0190_),
    .B(_0202_),
    .C(_0194_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4304_ (.I(net118),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4305_ (.I(_0189_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4306_ (.A1(_3326_),
    .A2(_0201_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4307_ (.I(_0193_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4308_ (.A1(_0203_),
    .A2(_0204_),
    .B(_0205_),
    .C(_0206_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4309_ (.I(net119),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4310_ (.A1(_3333_),
    .A2(_0201_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4311_ (.A1(_0207_),
    .A2(_0204_),
    .B(_0208_),
    .C(_0206_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4312_ (.I(net120),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4313_ (.A1(_3340_),
    .A2(_0201_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4314_ (.A1(_0209_),
    .A2(_0204_),
    .B(_0210_),
    .C(_0206_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4315_ (.I(net121),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4316_ (.I(_0200_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4317_ (.A1(_3348_),
    .A2(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4318_ (.A1(_0211_),
    .A2(_0204_),
    .B(_0213_),
    .C(_0206_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4319_ (.I(net122),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4320_ (.I(_0188_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4321_ (.I(_0215_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4322_ (.A1(_3356_),
    .A2(_0212_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4323_ (.I(_0193_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4324_ (.A1(_0214_),
    .A2(_0216_),
    .B(_0217_),
    .C(_0218_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4325_ (.I(net123),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4326_ (.A1(_3363_),
    .A2(_0212_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4327_ (.A1(_0219_),
    .A2(_0216_),
    .B(_0220_),
    .C(_0218_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4328_ (.I(net100),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4329_ (.A1(_3371_),
    .A2(_0212_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4330_ (.A1(_0221_),
    .A2(_0216_),
    .B(_0222_),
    .C(_0218_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4331_ (.I(net101),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4332_ (.I(_0200_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4333_ (.A1(_3379_),
    .A2(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4334_ (.A1(_0223_),
    .A2(_0216_),
    .B(_0225_),
    .C(_0218_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4335_ (.I(net102),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4336_ (.I(_0215_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4337_ (.A1(_3387_),
    .A2(_0224_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4338_ (.I(_0193_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4339_ (.A1(_0226_),
    .A2(_0227_),
    .B(_0228_),
    .C(_0229_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4340_ (.I(net103),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4341_ (.A1(_3393_),
    .A2(_0224_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4342_ (.A1(_0230_),
    .A2(_0227_),
    .B(_0231_),
    .C(_0229_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4343_ (.I(net104),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4344_ (.A1(_3401_),
    .A2(_0224_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4345_ (.A1(_0232_),
    .A2(_0227_),
    .B(_0233_),
    .C(_0229_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4346_ (.I(net105),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4347_ (.I(_0200_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4348_ (.A1(_3410_),
    .A2(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4349_ (.A1(_0234_),
    .A2(_0227_),
    .B(_0236_),
    .C(_0229_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4350_ (.I(net106),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4351_ (.I(_0215_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4352_ (.A1(_3417_),
    .A2(_0235_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4353_ (.I(net126),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4354_ (.I(_0240_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4355_ (.A1(_0237_),
    .A2(_0238_),
    .B(_0239_),
    .C(_0241_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4356_ (.I(net107),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4357_ (.A1(_3427_),
    .A2(_0235_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4358_ (.A1(_0242_),
    .A2(_0238_),
    .B(_0243_),
    .C(_0241_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4359_ (.I(net108),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4360_ (.A1(_3435_),
    .A2(_0235_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4361_ (.A1(_0244_),
    .A2(_0238_),
    .B(_0245_),
    .C(_0241_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4362_ (.I(net109),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4363_ (.I(_0188_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4364_ (.A1(_3444_),
    .A2(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4365_ (.A1(_0246_),
    .A2(_0238_),
    .B(_0248_),
    .C(_0241_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4366_ (.I(net111),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4367_ (.I(_0215_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4368_ (.A1(_3452_),
    .A2(_0247_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4369_ (.I(_0240_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4370_ (.A1(_0249_),
    .A2(_0250_),
    .B(_0251_),
    .C(_0252_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4371_ (.I(net112),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4372_ (.A1(_3461_),
    .A2(_0247_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4373_ (.A1(_0253_),
    .A2(_0250_),
    .B(_0254_),
    .C(_0252_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4374_ (.I(net113),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4375_ (.A1(_3469_),
    .A2(_0247_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4376_ (.A1(_0255_),
    .A2(_0250_),
    .B(_0256_),
    .C(_0252_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4377_ (.I(net114),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4378_ (.A1(_3475_),
    .A2(_0189_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4379_ (.A1(_0257_),
    .A2(_0250_),
    .B(_0258_),
    .C(_0252_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4380_ (.I(net115),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4381_ (.A1(_3483_),
    .A2(_0189_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4382_ (.I(_0240_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4383_ (.A1(_0259_),
    .A2(_0191_),
    .B(_0260_),
    .C(_0261_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4384_ (.I(_0163_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4385_ (.I(\dspArea_regB[0] ),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4386_ (.I(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4387_ (.I(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4388_ (.I(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4389_ (.I(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4390_ (.A1(_3283_),
    .A2(_3275_),
    .A3(_3279_),
    .A4(_0186_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4391_ (.I(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4392_ (.I0(_0267_),
    .I1(net99),
    .S(_0269_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4393_ (.A1(_0262_),
    .A2(_0270_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4394_ (.I(\dspArea_regB[1] ),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4395_ (.I(_0271_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4396_ (.I(_0272_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4397_ (.I(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4398_ (.I0(_0274_),
    .I1(net110),
    .S(_0269_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4399_ (.A1(_0262_),
    .A2(_0275_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4400_ (.I(\dspArea_regB[2] ),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4401_ (.I(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4402_ (.I(_0277_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4403_ (.I(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4404_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4405_ (.I0(_0280_),
    .I1(net116),
    .S(_0269_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4406_ (.A1(_0262_),
    .A2(_0281_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4407_ (.I(\dspArea_regB[3] ),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4408_ (.I(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4409_ (.I(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4410_ (.I(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4412_ (.I0(_0286_),
    .I1(net117),
    .S(_0269_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4413_ (.A1(_0262_),
    .A2(_0287_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4414_ (.I(_0163_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4415_ (.I(\dspArea_regB[4] ),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4416_ (.I(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4417_ (.I(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4418_ (.I(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4419_ (.I(_0268_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4420_ (.I0(_0292_),
    .I1(net118),
    .S(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4421_ (.A1(_0288_),
    .A2(_0294_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4422_ (.I(\dspArea_regB[5] ),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4423_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4424_ (.I(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4425_ (.I(_0297_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4426_ (.I0(_0298_),
    .I1(net119),
    .S(_0293_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4427_ (.A1(_0288_),
    .A2(_0299_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4428_ (.I(\dspArea_regB[6] ),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4429_ (.I(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4430_ (.I(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4431_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4432_ (.I0(_0303_),
    .I1(net120),
    .S(_0293_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4433_ (.A1(_0288_),
    .A2(_0304_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4434_ (.I(\dspArea_regB[7] ),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4435_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4436_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4437_ (.I(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4438_ (.I(_0308_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4439_ (.I0(_0309_),
    .I1(net121),
    .S(_0293_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4440_ (.A1(_0288_),
    .A2(_0310_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_0163_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4442_ (.I(\dspArea_regB[8] ),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4444_ (.I(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4445_ (.I(_0314_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4446_ (.I(_0268_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4447_ (.I0(_0315_),
    .I1(net122),
    .S(_0316_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4448_ (.A1(_0311_),
    .A2(_0317_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4449_ (.I(\dspArea_regB[9] ),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4450_ (.I(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4451_ (.I(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4452_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4453_ (.I(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4454_ (.I(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4455_ (.I0(_0323_),
    .I1(net123),
    .S(_0316_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4456_ (.A1(_0311_),
    .A2(_0324_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4457_ (.I(\dspArea_regB[10] ),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4458_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4459_ (.I(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4460_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4461_ (.I0(_0328_),
    .I1(net100),
    .S(_0316_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4462_ (.A1(_0311_),
    .A2(_0329_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4463_ (.I(\dspArea_regB[11] ),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4464_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4465_ (.I(_0331_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4466_ (.I(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4467_ (.I(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4468_ (.I(_0334_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4469_ (.I0(_0335_),
    .I1(net101),
    .S(_0316_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4470_ (.A1(_0311_),
    .A2(_0336_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4471_ (.I(_3487_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4472_ (.I(_0337_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4473_ (.I(\dspArea_regB[12] ),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4474_ (.I(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4475_ (.I(_0340_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4476_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4477_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4478_ (.I(_0268_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4479_ (.I0(_0343_),
    .I1(net102),
    .S(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4480_ (.A1(_0338_),
    .A2(_0345_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4481_ (.I(\dspArea_regB[13] ),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4482_ (.I(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4483_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4485_ (.I(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4486_ (.I0(_0350_),
    .I1(net103),
    .S(_0344_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4487_ (.A1(_0338_),
    .A2(_0351_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4488_ (.I(\dspArea_regB[14] ),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4489_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4490_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4491_ (.I(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4492_ (.I(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4493_ (.I0(_0356_),
    .I1(net104),
    .S(_0344_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4494_ (.A1(_0338_),
    .A2(_0357_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(\dspArea_regB[15] ),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4496_ (.I(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4497_ (.I(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4498_ (.I(_0360_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4499_ (.I(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4500_ (.I0(_0362_),
    .I1(net105),
    .S(_0344_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4501_ (.A1(_0338_),
    .A2(_0363_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(_0337_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4503_ (.A1(_3274_),
    .A2(_3284_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4504_ (.I(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4505_ (.A1(net98),
    .A2(net159),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4506_ (.A1(net125),
    .A2(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4507_ (.A1(_3271_),
    .A2(_3286_),
    .A3(_0366_),
    .A4(_0368_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4508_ (.I(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4509_ (.A1(_0267_),
    .A2(_3294_),
    .A3(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4510_ (.A1(\dspArea_regP[0] ),
    .A2(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4511_ (.A1(_0364_),
    .A2(_0372_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4512_ (.A1(\dspArea_regP[0] ),
    .A2(_0267_),
    .A3(_3294_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4513_ (.A1(_0267_),
    .A2(_3301_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4514_ (.A1(\dspArea_regP[1] ),
    .A2(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4515_ (.A1(_0274_),
    .A2(_3293_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4516_ (.A1(_0375_),
    .A2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4517_ (.A1(_0373_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4518_ (.I(_0369_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4519_ (.I(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4520_ (.I0(\dspArea_regP[1] ),
    .I1(_0378_),
    .S(_0380_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4521_ (.A1(_0364_),
    .A2(_0381_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4522_ (.A1(_0373_),
    .A2(_0377_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4523_ (.A1(_0266_),
    .A2(_3307_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4524_ (.A1(\dspArea_regP[2] ),
    .A2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4525_ (.A1(_0274_),
    .A2(_3302_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4526_ (.A1(_0384_),
    .A2(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4527_ (.A1(\dspArea_regP[1] ),
    .A2(_0374_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4528_ (.A1(_0375_),
    .A2(_0376_),
    .B(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4529_ (.A1(_0386_),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4530_ (.I(_3291_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4531_ (.I(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4532_ (.A1(_0280_),
    .A2(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4533_ (.A1(_0389_),
    .A2(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4534_ (.A1(_0382_),
    .A2(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4535_ (.I(_0369_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4536_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4537_ (.I0(\dspArea_regP[2] ),
    .I1(_0394_),
    .S(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4538_ (.A1(_0364_),
    .A2(_0397_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4539_ (.A1(_0382_),
    .A2(_0393_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4540_ (.A1(_0274_),
    .A2(_3307_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4541_ (.I(_3314_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4542_ (.A1(_0266_),
    .A2(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4543_ (.A1(\dspArea_regP[3] ),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4544_ (.A1(_0399_),
    .A2(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4545_ (.A1(\dspArea_regP[2] ),
    .A2(_0383_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4546_ (.A1(_0384_),
    .A2(_0385_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4547_ (.A1(_0403_),
    .A2(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4548_ (.A1(_0280_),
    .A2(_3301_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4549_ (.A1(_0286_),
    .A2(_3293_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4550_ (.A1(_0285_),
    .A2(_3300_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4551_ (.A1(_0392_),
    .A2(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4552_ (.A1(_0407_),
    .A2(_0408_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4553_ (.A1(_0406_),
    .A2(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4554_ (.I(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4555_ (.I(_0386_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4556_ (.A1(_0414_),
    .A2(_0388_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4557_ (.A1(_0280_),
    .A2(_3293_),
    .A3(_0389_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4558_ (.A1(_0415_),
    .A2(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4559_ (.A1(_0413_),
    .A2(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4560_ (.A1(_0398_),
    .A2(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4561_ (.I0(\dspArea_regP[3] ),
    .I1(_0419_),
    .S(_0396_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4562_ (.A1(_0364_),
    .A2(_0420_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4563_ (.I(\dspArea_regP[4] ),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4564_ (.A1(_3288_),
    .A2(_0368_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4565_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4566_ (.I(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4567_ (.A1(_3287_),
    .A2(_0368_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4568_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4569_ (.A1(_0279_),
    .A2(_3305_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4570_ (.A1(_0409_),
    .A2(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4571_ (.A1(_0292_),
    .A2(_3292_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4572_ (.A1(_0428_),
    .A2(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4573_ (.I(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4574_ (.A1(_0273_),
    .A2(_0400_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4575_ (.I(_3321_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4576_ (.A1(_0266_),
    .A2(_0433_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4577_ (.A1(\dspArea_regP[4] ),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4578_ (.A1(_0432_),
    .A2(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4579_ (.A1(\dspArea_regP[3] ),
    .A2(_0401_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4580_ (.A1(_0399_),
    .A2(_0402_),
    .B(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4581_ (.A1(_0431_),
    .A2(_0436_),
    .A3(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4582_ (.A1(_0403_),
    .A2(_0405_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4583_ (.I(_0411_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4584_ (.A1(_0406_),
    .A2(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4585_ (.A1(_0440_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4586_ (.A1(_0410_),
    .A2(_0439_),
    .A3(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4587_ (.A1(_0413_),
    .A2(_0417_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4588_ (.A1(_0398_),
    .A2(_0418_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4589_ (.A1(_0445_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4590_ (.A1(_0444_),
    .A2(_0447_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4591_ (.A1(_0444_),
    .A2(_0447_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4592_ (.A1(_0426_),
    .A2(_0448_),
    .A3(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4593_ (.A1(_0421_),
    .A2(_0424_),
    .B(_0450_),
    .C(_0261_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4594_ (.I(_0426_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4595_ (.A1(_0446_),
    .A2(_0444_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4596_ (.A1(_0445_),
    .A2(_0444_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4597_ (.A1(_0286_),
    .A2(_3307_),
    .A3(_0407_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4598_ (.A1(_0292_),
    .A2(_3292_),
    .A3(_0428_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4599_ (.A1(_0454_),
    .A2(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4600_ (.A1(_0298_),
    .A2(_3290_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4601_ (.A1(_0456_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4602_ (.I(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4603_ (.I(_0290_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4604_ (.I(_3299_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4605_ (.I(_0461_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4606_ (.A1(_0460_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4607_ (.I(_0282_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4608_ (.I(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4609_ (.I(_3304_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4610_ (.A1(_0465_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4611_ (.I(\dspArea_regB[2] ),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4613_ (.I(_0469_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4614_ (.A1(_0470_),
    .A2(_3314_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4615_ (.A1(_0467_),
    .A2(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4616_ (.A1(_0463_),
    .A2(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4617_ (.I(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4618_ (.A1(_0273_),
    .A2(_0433_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4619_ (.I(_0263_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4620_ (.I(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4621_ (.I(_3328_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4622_ (.A1(_0477_),
    .A2(_0478_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4623_ (.A1(\dspArea_regP[5] ),
    .A2(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4624_ (.A1(_0475_),
    .A2(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4625_ (.A1(\dspArea_regP[4] ),
    .A2(_0434_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4626_ (.A1(_0432_),
    .A2(_0435_),
    .B(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4627_ (.A1(_0474_),
    .A2(_0481_),
    .A3(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4628_ (.A1(_0436_),
    .A2(_0438_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4629_ (.A1(_0436_),
    .A2(_0438_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4630_ (.A1(_0431_),
    .A2(_0485_),
    .B(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4631_ (.A1(_0459_),
    .A2(_0484_),
    .A3(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4632_ (.A1(_0440_),
    .A2(_0442_),
    .A3(_0439_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4633_ (.A1(_0440_),
    .A2(_0442_),
    .B(_0439_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4634_ (.A1(_0410_),
    .A2(_0489_),
    .B(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4635_ (.A1(_0488_),
    .A2(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4636_ (.A1(_0453_),
    .A2(_0492_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4637_ (.A1(_0452_),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4638_ (.I(_0425_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4639_ (.A1(\dspArea_regP[5] ),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4640_ (.A1(_0451_),
    .A2(_0494_),
    .B(_0496_),
    .C(_0261_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(_0337_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4642_ (.A1(_0452_),
    .A2(_0493_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4643_ (.A1(_0454_),
    .A2(_0455_),
    .B(_0457_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4644_ (.A1(_0286_),
    .A2(_0400_),
    .A3(_0427_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4645_ (.I(_3300_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4646_ (.A1(_0292_),
    .A2(_0501_),
    .A3(_0472_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4647_ (.A1(_0500_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4648_ (.A1(_0298_),
    .A2(_3300_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4649_ (.A1(_0303_),
    .A2(_3291_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4650_ (.A1(_0504_),
    .A2(_0505_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4651_ (.I(\dspArea_regB[6] ),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4652_ (.A1(_0507_),
    .A2(\dspArea_regA[1] ),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4653_ (.A1(_0457_),
    .A2(_0508_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4654_ (.A1(_0506_),
    .A2(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4655_ (.A1(_0503_),
    .A2(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4656_ (.I(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4657_ (.A1(_0290_),
    .A2(_0466_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4658_ (.I(\dspArea_regB[3] ),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4659_ (.I(_0514_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4660_ (.A1(_0515_),
    .A2(_3312_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4661_ (.A1(_0468_),
    .A2(_3321_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4662_ (.A1(_0516_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4663_ (.A1(_0513_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4664_ (.I(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4665_ (.I(_3329_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4666_ (.A1(\dspArea_regP[5] ),
    .A2(_0265_),
    .A3(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4667_ (.I(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4668_ (.A1(_0475_),
    .A2(_0480_),
    .B(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4669_ (.A1(_0273_),
    .A2(_3331_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4670_ (.A1(_0265_),
    .A2(_3337_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4671_ (.A1(\dspArea_regP[6] ),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4672_ (.A1(_0525_),
    .A2(_0527_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4673_ (.A1(_0520_),
    .A2(_0524_),
    .A3(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4674_ (.A1(_0481_),
    .A2(_0483_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4675_ (.A1(_0481_),
    .A2(_0483_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4676_ (.A1(_0474_),
    .A2(_0530_),
    .B(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4677_ (.A1(_0529_),
    .A2(_0532_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4678_ (.A1(_0512_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4679_ (.A1(_0484_),
    .A2(_0487_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4680_ (.A1(_0484_),
    .A2(_0487_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4681_ (.A1(_0459_),
    .A2(_0535_),
    .B(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4682_ (.A1(_0499_),
    .A2(_0534_),
    .A3(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4683_ (.A1(_0488_),
    .A2(_0491_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4684_ (.A1(_0453_),
    .A2(_0492_),
    .B(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4685_ (.A1(_0538_),
    .A2(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4686_ (.A1(_0498_),
    .A2(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4687_ (.I0(\dspArea_regP[6] ),
    .I1(_0542_),
    .S(_0396_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4688_ (.A1(_0497_),
    .A2(_0543_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4689_ (.A1(_0498_),
    .A2(_0541_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4690_ (.A1(_0488_),
    .A2(_0491_),
    .A3(_0538_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4691_ (.A1(_0503_),
    .A2(_0510_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4692_ (.I(_0283_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4693_ (.A1(_0547_),
    .A2(_3324_),
    .A3(_0471_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4694_ (.A1(_0291_),
    .A2(_3305_),
    .A3(_0518_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4695_ (.A1(_0548_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4696_ (.I(_0305_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4697_ (.I(\dspArea_regA[0] ),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4698_ (.A1(_0551_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4699_ (.I(\dspArea_regB[5] ),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4700_ (.I(\dspArea_regA[2] ),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4701_ (.A1(_0554_),
    .A2(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4702_ (.A1(_0508_),
    .A2(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4703_ (.A1(_0553_),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4704_ (.A1(_0550_),
    .A2(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4705_ (.A1(_0509_),
    .A2(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4706_ (.I(_0289_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4707_ (.I(_0561_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4708_ (.A1(_0562_),
    .A2(_3315_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4709_ (.I(_0282_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4710_ (.A1(_0564_),
    .A2(_3322_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4711_ (.A1(_0469_),
    .A2(_3329_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4712_ (.A1(_0565_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4713_ (.A1(_0563_),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4714_ (.I(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4715_ (.I(_0272_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4716_ (.A1(_0570_),
    .A2(_3338_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4717_ (.A1(_0477_),
    .A2(_3344_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4718_ (.A1(\dspArea_regP[7] ),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4719_ (.A1(_0571_),
    .A2(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4720_ (.A1(\dspArea_regP[6] ),
    .A2(_0526_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4721_ (.A1(_0525_),
    .A2(_0527_),
    .B(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4722_ (.A1(_0569_),
    .A2(_0574_),
    .A3(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4723_ (.A1(_0524_),
    .A2(_0528_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4724_ (.A1(_0524_),
    .A2(_0528_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4725_ (.A1(_0520_),
    .A2(_0578_),
    .B(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4726_ (.A1(_0560_),
    .A2(_0577_),
    .A3(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4727_ (.A1(_0529_),
    .A2(_0532_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4728_ (.A1(_0529_),
    .A2(_0532_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4729_ (.A1(_0512_),
    .A2(_0582_),
    .B(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4730_ (.A1(_0581_),
    .A2(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4731_ (.A1(_0546_),
    .A2(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4732_ (.A1(_0534_),
    .A2(_0537_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4733_ (.A1(_0534_),
    .A2(_0537_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4734_ (.A1(_0499_),
    .A2(_0587_),
    .B(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4735_ (.A1(_0545_),
    .A2(_0586_),
    .A3(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4736_ (.A1(_0453_),
    .A2(_0492_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4737_ (.A1(_0591_),
    .A2(_0538_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4738_ (.A1(_0544_),
    .A2(_0590_),
    .A3(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4739_ (.I0(\dspArea_regP[7] ),
    .I1(_0593_),
    .S(_0396_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4740_ (.A1(_0497_),
    .A2(_0594_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4741_ (.A1(_0590_),
    .A2(_0592_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4742_ (.A1(_0590_),
    .A2(_0592_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4743_ (.A1(_0544_),
    .A2(_0595_),
    .B(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4744_ (.I(_0550_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4745_ (.A1(_0598_),
    .A2(_0558_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4746_ (.A1(_0509_),
    .A2(_0559_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4747_ (.A1(_0599_),
    .A2(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4748_ (.A1(_0315_),
    .A2(_3291_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4749_ (.A1(_0601_),
    .A2(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4750_ (.I(_0300_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4751_ (.A1(_0604_),
    .A2(_0555_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4752_ (.A1(_0504_),
    .A2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4753_ (.I(_0551_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4754_ (.I(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4755_ (.A1(_0608_),
    .A2(_3290_),
    .A3(_0557_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4756_ (.A1(_0606_),
    .A2(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4757_ (.A1(_0547_),
    .A2(_0521_),
    .A3(_0517_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4758_ (.A1(_0291_),
    .A2(_3315_),
    .A3(_0567_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4759_ (.A1(_0611_),
    .A2(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4760_ (.I(\dspArea_regB[7] ),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4761_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4762_ (.A1(_0615_),
    .A2(_0461_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4763_ (.A1(_0554_),
    .A2(_3313_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4764_ (.A1(_0605_),
    .A2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4765_ (.A1(_0616_),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4766_ (.A1(_0613_),
    .A2(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4767_ (.A1(_0610_),
    .A2(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4768_ (.I(\dspArea_regB[4] ),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4769_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4770_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4771_ (.A1(_0624_),
    .A2(_3323_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4772_ (.A1(_0515_),
    .A2(_3329_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4773_ (.A1(_0277_),
    .A2(_3335_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4774_ (.A1(_0626_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4775_ (.A1(_0625_),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4776_ (.I(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4777_ (.I(_3345_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4778_ (.A1(_0272_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4779_ (.A1(_0264_),
    .A2(_3352_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4780_ (.A1(\dspArea_regP[8] ),
    .A2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4781_ (.A1(_0632_),
    .A2(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4782_ (.A1(\dspArea_regP[7] ),
    .A2(_0572_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4783_ (.A1(_0571_),
    .A2(_0573_),
    .B(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4784_ (.A1(_0630_),
    .A2(_0635_),
    .A3(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4785_ (.A1(_0574_),
    .A2(_0576_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4786_ (.A1(_0574_),
    .A2(_0576_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4787_ (.A1(_0569_),
    .A2(_0639_),
    .B(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4788_ (.A1(_0638_),
    .A2(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4789_ (.A1(_0621_),
    .A2(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4790_ (.A1(_0577_),
    .A2(_0580_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4791_ (.A1(_0577_),
    .A2(_0580_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4792_ (.A1(_0560_),
    .A2(_0644_),
    .B(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4793_ (.A1(_0643_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4794_ (.A1(_0603_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4795_ (.A1(_0511_),
    .A2(_0533_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4796_ (.A1(_0583_),
    .A2(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4797_ (.A1(_0503_),
    .A2(_0510_),
    .A3(_0585_),
    .B1(_0650_),
    .B2(_0581_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4798_ (.A1(_0648_),
    .A2(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4799_ (.A1(_0586_),
    .A2(_0589_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4800_ (.A1(_0586_),
    .A2(_0589_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4801_ (.A1(_0545_),
    .A2(_0653_),
    .B(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4802_ (.A1(_0652_),
    .A2(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4803_ (.A1(_0597_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4804_ (.A1(\dspArea_regP[8] ),
    .A2(_0495_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4805_ (.A1(_0451_),
    .A2(_0657_),
    .B(_0658_),
    .C(_0261_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4806_ (.A1(_0597_),
    .A2(_0656_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4807_ (.A1(_0545_),
    .A2(_0653_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4808_ (.A1(_0660_),
    .A2(_0652_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4809_ (.A1(_0601_),
    .A2(_0602_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4810_ (.I(_0613_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4811_ (.A1(_0663_),
    .A2(_0619_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4812_ (.A1(_0610_),
    .A2(_0620_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4813_ (.A1(_0664_),
    .A2(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4814_ (.A1(_0315_),
    .A2(_0462_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4815_ (.A1(_0323_),
    .A2(_0391_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4816_ (.A1(_0666_),
    .A2(_0667_),
    .A3(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4817_ (.I(_3313_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4818_ (.A1(_0301_),
    .A2(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4819_ (.A1(_0556_),
    .A2(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4820_ (.A1(_0309_),
    .A2(_0501_),
    .A3(_0618_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4821_ (.A1(_0672_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4822_ (.I(_0284_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4823_ (.A1(_0675_),
    .A2(_3338_),
    .A3(_0566_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4824_ (.I(_0622_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4825_ (.I(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4826_ (.A1(_0678_),
    .A2(_3324_),
    .A3(_0628_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4827_ (.A1(_0676_),
    .A2(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4828_ (.A1(_0607_),
    .A2(_3305_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4829_ (.A1(_0297_),
    .A2(_3322_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4830_ (.A1(_0671_),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4831_ (.A1(_0681_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4832_ (.A1(_0680_),
    .A2(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4833_ (.A1(_0674_),
    .A2(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4834_ (.A1(_0677_),
    .A2(_0521_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4835_ (.A1(_0464_),
    .A2(_3336_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4836_ (.I(_3343_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4837_ (.A1(_0277_),
    .A2(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4838_ (.A1(_0688_),
    .A2(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4839_ (.A1(_0687_),
    .A2(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4840_ (.I(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4841_ (.I(\dspArea_regB[1] ),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4842_ (.I(_3352_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4843_ (.A1(_0694_),
    .A2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4844_ (.I(_0263_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4845_ (.A1(_0697_),
    .A2(\dspArea_regA[9] ),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4846_ (.A1(\dspArea_regP[9] ),
    .A2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4847_ (.A1(_0696_),
    .A2(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4848_ (.A1(\dspArea_regP[8] ),
    .A2(_0633_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4849_ (.A1(_0632_),
    .A2(_0634_),
    .B(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4850_ (.A1(_0700_),
    .A2(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4851_ (.A1(_0693_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4852_ (.A1(_0635_),
    .A2(_0637_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4853_ (.A1(_0635_),
    .A2(_0637_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4854_ (.A1(_0630_),
    .A2(_0705_),
    .B(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4855_ (.A1(_0704_),
    .A2(_0707_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4856_ (.A1(_0686_),
    .A2(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4857_ (.A1(_0638_),
    .A2(_0641_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4858_ (.A1(_0621_),
    .A2(_0642_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4859_ (.A1(_0710_),
    .A2(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4860_ (.A1(_0669_),
    .A2(_0709_),
    .A3(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4861_ (.A1(_0643_),
    .A2(_0646_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4862_ (.A1(_0603_),
    .A2(_0647_),
    .B(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4863_ (.A1(_0713_),
    .A2(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4864_ (.A1(_0662_),
    .A2(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4865_ (.A1(_0603_),
    .A2(_0647_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4866_ (.A1(_0718_),
    .A2(_0651_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4867_ (.A1(_0654_),
    .A2(_0652_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4868_ (.A1(_0719_),
    .A2(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4869_ (.A1(_0717_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4870_ (.A1(_0659_),
    .A2(_0661_),
    .B(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4871_ (.A1(_0659_),
    .A2(_0661_),
    .A3(_0722_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4872_ (.A1(_0723_),
    .A2(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4873_ (.I(_0395_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4874_ (.I0(\dspArea_regP[9] ),
    .I1(_0725_),
    .S(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4875_ (.A1(_0497_),
    .A2(_0727_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4876_ (.A1(_0717_),
    .A2(_0720_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4877_ (.A1(_0723_),
    .A2(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4878_ (.A1(_0719_),
    .A2(_0717_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4879_ (.A1(_0713_),
    .A2(_0715_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4880_ (.A1(_0662_),
    .A2(_0716_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4881_ (.A1(_0731_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4882_ (.A1(_0667_),
    .A2(_0668_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4883_ (.I(\dspArea_regB[9] ),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4884_ (.I(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4885_ (.I(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4886_ (.A1(_0737_),
    .A2(_3299_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4887_ (.A1(_0602_),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4888_ (.A1(_0666_),
    .A2(_0734_),
    .A3(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4889_ (.I(_0680_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4890_ (.A1(_0741_),
    .A2(_0684_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4891_ (.A1(_0674_),
    .A2(_0685_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4892_ (.A1(_0742_),
    .A2(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4893_ (.A1(_0314_),
    .A2(_3304_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4894_ (.A1(_0738_),
    .A2(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4895_ (.I(\dspArea_regB[10] ),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4896_ (.I(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4897_ (.A1(_0748_),
    .A2(_3290_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4898_ (.A1(_0746_),
    .A2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4899_ (.A1(_0739_),
    .A2(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4900_ (.A1(_0744_),
    .A2(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4901_ (.A1(_0303_),
    .A2(_3325_),
    .A3(_0617_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4902_ (.A1(_0309_),
    .A2(_3306_),
    .A3(_0683_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4903_ (.A1(_0753_),
    .A2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4904_ (.A1(_0564_),
    .A2(_3344_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4905_ (.A1(_0627_),
    .A2(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4906_ (.A1(_0678_),
    .A2(_3331_),
    .A3(_0691_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4907_ (.A1(_0757_),
    .A2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4908_ (.I(_0615_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4909_ (.A1(_0760_),
    .A2(_3315_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4910_ (.A1(_0301_),
    .A2(_3323_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4911_ (.A1(_0297_),
    .A2(_0478_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4912_ (.A1(_0762_),
    .A2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4913_ (.A1(_0761_),
    .A2(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4914_ (.A1(_0759_),
    .A2(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4915_ (.A1(_0755_),
    .A2(_0766_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4916_ (.I(\dspArea_regB[4] ),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4917_ (.I(_3336_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4918_ (.A1(_0768_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4919_ (.A1(_0470_),
    .A2(_3353_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4920_ (.A1(_0756_),
    .A2(_0770_),
    .A3(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4921_ (.I(_3359_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4922_ (.A1(_0272_),
    .A2(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4923_ (.A1(_0264_),
    .A2(_3366_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4924_ (.A1(\dspArea_regP[10] ),
    .A2(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4925_ (.A1(_0774_),
    .A2(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4926_ (.A1(\dspArea_regP[9] ),
    .A2(_0698_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4927_ (.A1(_0696_),
    .A2(_0699_),
    .B(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4928_ (.A1(_0772_),
    .A2(_0777_),
    .A3(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4929_ (.A1(_0700_),
    .A2(_0702_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4930_ (.A1(_0700_),
    .A2(_0702_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4931_ (.A1(_0693_),
    .A2(_0781_),
    .B(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4932_ (.A1(_0780_),
    .A2(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4933_ (.A1(_0767_),
    .A2(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4934_ (.A1(_0704_),
    .A2(_0707_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4935_ (.A1(_0686_),
    .A2(_0708_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4936_ (.A1(_0786_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4937_ (.A1(_0752_),
    .A2(_0785_),
    .A3(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4938_ (.A1(_0710_),
    .A2(_0711_),
    .A3(_0709_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4939_ (.A1(_0710_),
    .A2(_0711_),
    .B(_0709_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4940_ (.A1(_0669_),
    .A2(_0790_),
    .B(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4941_ (.A1(_0789_),
    .A2(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4942_ (.A1(_0740_),
    .A2(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4943_ (.A1(_0730_),
    .A2(_0733_),
    .A3(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4944_ (.I(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4945_ (.A1(_0729_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4946_ (.I0(\dspArea_regP[10] ),
    .I1(_0797_),
    .S(_0726_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4947_ (.A1(_0497_),
    .A2(_0798_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4948_ (.I(_0370_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4949_ (.A1(\dspArea_regP[11] ),
    .A2(_0799_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4950_ (.A1(_0731_),
    .A2(_0732_),
    .A3(_0794_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4951_ (.A1(_0731_),
    .A2(_0732_),
    .B(_0794_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4952_ (.A1(_0730_),
    .A2(_0801_),
    .A3(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4953_ (.A1(_0729_),
    .A2(_0795_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4954_ (.A1(_0803_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4955_ (.I(_0802_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4956_ (.A1(_0744_),
    .A2(_0751_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4957_ (.I(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4958_ (.A1(_0739_),
    .A2(_0750_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4959_ (.I(_0759_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4960_ (.A1(_0810_),
    .A2(_0765_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4961_ (.A1(_0755_),
    .A2(_0766_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4962_ (.A1(_0811_),
    .A2(_0812_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4963_ (.A1(_0327_),
    .A2(_0462_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4964_ (.I(_0318_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4965_ (.A1(_0815_),
    .A2(\dspArea_regA[2] ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4966_ (.A1(_0313_),
    .A2(_3312_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4967_ (.A1(_0816_),
    .A2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4968_ (.A1(_0814_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4969_ (.A1(_0667_),
    .A2(_0816_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4970_ (.A1(_0748_),
    .A2(_0552_),
    .A3(_0746_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4971_ (.A1(_0820_),
    .A2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4972_ (.A1(_0819_),
    .A2(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4973_ (.A1(_0335_),
    .A2(_3292_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4974_ (.A1(_0823_),
    .A2(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4975_ (.I(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4976_ (.A1(_0809_),
    .A2(_0813_),
    .A3(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4977_ (.I(_0301_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4978_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4979_ (.A1(_0829_),
    .A2(_3331_),
    .A3(_0682_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4980_ (.A1(_0608_),
    .A2(_0400_),
    .A3(_0764_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4981_ (.A1(_0830_),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4982_ (.A1(_0756_),
    .A2(_0771_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4983_ (.I(_0695_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4984_ (.A1(_0465_),
    .A2(_0470_),
    .A3(_0834_),
    .A4(_0631_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4985_ (.I(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4986_ (.A1(_0770_),
    .A2(_0833_),
    .B(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4987_ (.A1(_0306_),
    .A2(_3323_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4988_ (.I(_0300_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4989_ (.A1(_0839_),
    .A2(_0478_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4990_ (.A1(_0296_),
    .A2(_3335_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4991_ (.A1(_0840_),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4992_ (.A1(_0838_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4993_ (.A1(_0837_),
    .A2(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4994_ (.A1(_0832_),
    .A2(_0844_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4995_ (.A1(_0283_),
    .A2(_3353_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4996_ (.A1(_0561_),
    .A2(_3345_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4997_ (.A1(_0279_),
    .A2(_3360_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4998_ (.A1(_0846_),
    .A2(_0847_),
    .A3(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4999_ (.I(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5000_ (.A1(_0570_),
    .A2(_3368_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5001_ (.A1(_0477_),
    .A2(_3375_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5002_ (.A1(\dspArea_regP[11] ),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5003_ (.A1(_0851_),
    .A2(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5004_ (.A1(\dspArea_regP[10] ),
    .A2(_0775_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5005_ (.A1(_0774_),
    .A2(_0776_),
    .B(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5006_ (.A1(_0850_),
    .A2(_0854_),
    .A3(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5007_ (.I(_0772_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5008_ (.A1(_0777_),
    .A2(_0779_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5009_ (.A1(_0777_),
    .A2(_0779_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5010_ (.A1(_0858_),
    .A2(_0859_),
    .B(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5011_ (.A1(_0857_),
    .A2(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5012_ (.A1(_0845_),
    .A2(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5013_ (.A1(_0692_),
    .A2(_0703_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5014_ (.A1(_0782_),
    .A2(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5015_ (.A1(_0780_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5016_ (.A1(_0767_),
    .A2(_0784_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5017_ (.A1(_0866_),
    .A2(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5018_ (.A1(_0827_),
    .A2(_0863_),
    .A3(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5019_ (.A1(_0786_),
    .A2(_0787_),
    .A3(_0785_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5020_ (.A1(_0786_),
    .A2(_0787_),
    .B(_0785_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5021_ (.A1(_0752_),
    .A2(_0870_),
    .B(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5022_ (.A1(_0808_),
    .A2(_0869_),
    .A3(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5023_ (.A1(_0789_),
    .A2(_0792_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5024_ (.A1(_0740_),
    .A2(_0793_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5025_ (.A1(_0874_),
    .A2(_0875_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5026_ (.A1(_0873_),
    .A2(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5027_ (.A1(_0806_),
    .A2(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5028_ (.A1(_0805_),
    .A2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5029_ (.A1(_0805_),
    .A2(_0878_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5030_ (.A1(_0423_),
    .A2(_0879_),
    .A3(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5031_ (.A1(_3681_),
    .A2(_0800_),
    .A3(_0881_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5032_ (.I(_0337_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5033_ (.A1(_0597_),
    .A2(_0656_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5034_ (.A1(_0660_),
    .A2(_0652_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5035_ (.I(_0717_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5036_ (.A1(_0885_),
    .A2(_0721_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5037_ (.A1(_0885_),
    .A2(_0721_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5038_ (.A1(_0883_),
    .A2(_0884_),
    .B(_0886_),
    .C(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5039_ (.I(_0728_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5040_ (.A1(_0806_),
    .A2(_0877_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5041_ (.A1(_0806_),
    .A2(_0877_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5042_ (.A1(_0888_),
    .A2(_0889_),
    .B1(_0890_),
    .B2(_0891_),
    .C(_0795_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5043_ (.I(_0877_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5044_ (.A1(_0806_),
    .A2(_0803_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5045_ (.A1(_0893_),
    .A2(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5046_ (.A1(_0892_),
    .A2(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5047_ (.I(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5048_ (.I(_0873_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5049_ (.A1(_0869_),
    .A2(_0872_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5050_ (.A1(_0869_),
    .A2(_0872_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5051_ (.A1(_0808_),
    .A2(_0899_),
    .B(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5052_ (.A1(_0813_),
    .A2(_0826_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5053_ (.A1(_0813_),
    .A2(_0826_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5054_ (.A1(_0809_),
    .A2(_0903_),
    .A3(_0902_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5055_ (.A1(_0902_),
    .A2(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5056_ (.I(_0822_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5057_ (.A1(_0819_),
    .A2(_0906_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5058_ (.A1(_0335_),
    .A2(_0390_),
    .A3(_0823_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5059_ (.A1(_0907_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5060_ (.I(_0843_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5061_ (.A1(_0837_),
    .A2(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5062_ (.A1(_0832_),
    .A2(_0844_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5063_ (.A1(_0911_),
    .A2(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5064_ (.A1(_0333_),
    .A2(_0462_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5065_ (.I(_0341_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5066_ (.A1(_0915_),
    .A2(_0552_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5067_ (.A1(_0914_),
    .A2(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5068_ (.A1(_0747_),
    .A2(_0466_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5069_ (.A1(_0815_),
    .A2(_3312_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5070_ (.I(\dspArea_regA[4] ),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5071_ (.A1(_0313_),
    .A2(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5072_ (.A1(_0919_),
    .A2(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5073_ (.A1(_0918_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5074_ (.I(_0320_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5075_ (.A1(_0924_),
    .A2(_3314_),
    .A3(_0745_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5076_ (.I(\dspArea_regB[10] ),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5077_ (.I(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5078_ (.I(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5079_ (.A1(_0928_),
    .A2(_0461_),
    .A3(_0818_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5080_ (.A1(_0925_),
    .A2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5081_ (.A1(_0923_),
    .A2(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5082_ (.A1(_0917_),
    .A2(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5083_ (.A1(_0913_),
    .A2(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5084_ (.A1(_0909_),
    .A2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5085_ (.A1(_0303_),
    .A2(_3339_),
    .A3(_0763_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5086_ (.A1(_0838_),
    .A2(_0842_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5087_ (.A1(_0935_),
    .A2(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5088_ (.A1(_0846_),
    .A2(_0848_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _5089_ (.A1(_0465_),
    .A2(_0470_),
    .A3(_0773_),
    .A4(_0834_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5090_ (.I(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5091_ (.A1(_0847_),
    .A2(_0938_),
    .B(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5092_ (.A1(_0614_),
    .A2(_3330_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5093_ (.A1(_0507_),
    .A2(_3336_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5094_ (.A1(_0296_),
    .A2(_0689_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5095_ (.A1(_0943_),
    .A2(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5096_ (.A1(_0942_),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5097_ (.A1(_0941_),
    .A2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5098_ (.A1(_0937_),
    .A2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5099_ (.I(\dspArea_regA[9] ),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5100_ (.A1(_0564_),
    .A2(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5101_ (.A1(_0768_),
    .A2(_0695_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5102_ (.A1(_0278_),
    .A2(_3367_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5103_ (.A1(_0950_),
    .A2(_0951_),
    .A3(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5104_ (.I(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5105_ (.I(\dspArea_regA[11] ),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5106_ (.I(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5107_ (.A1(_0570_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5108_ (.I(\dspArea_regA[12] ),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5109_ (.I(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5110_ (.A1(_0477_),
    .A2(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5111_ (.A1(\dspArea_regP[12] ),
    .A2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5112_ (.A1(_0957_),
    .A2(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5113_ (.A1(\dspArea_regP[11] ),
    .A2(_0852_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5114_ (.A1(_0851_),
    .A2(_0853_),
    .B(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5115_ (.A1(_0954_),
    .A2(_0962_),
    .A3(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5116_ (.A1(_0854_),
    .A2(_0856_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5117_ (.A1(_0854_),
    .A2(_0856_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5118_ (.A1(_0850_),
    .A2(_0966_),
    .B(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5119_ (.A1(_0965_),
    .A2(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5120_ (.A1(_0948_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5121_ (.A1(_0857_),
    .A2(_0861_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5122_ (.A1(_0845_),
    .A2(_0862_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5123_ (.A1(_0971_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5124_ (.A1(_0934_),
    .A2(_0970_),
    .A3(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5125_ (.A1(_0866_),
    .A2(_0867_),
    .A3(_0863_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5126_ (.A1(_0866_),
    .A2(_0867_),
    .B(_0863_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5127_ (.A1(_0827_),
    .A2(_0975_),
    .B(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5128_ (.A1(_0974_),
    .A2(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5129_ (.A1(_0901_),
    .A2(_0905_),
    .A3(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5130_ (.A1(_0898_),
    .A2(_0876_),
    .B(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5131_ (.A1(_0898_),
    .A2(_0876_),
    .A3(_0979_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5132_ (.A1(_0980_),
    .A2(_0981_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5133_ (.A1(_0897_),
    .A2(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5134_ (.I0(\dspArea_regP[12] ),
    .I1(_0983_),
    .S(_0726_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5135_ (.A1(_0882_),
    .A2(_0984_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5136_ (.A1(_3271_),
    .A2(_3277_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _5137_ (.A1(net125),
    .A2(_3276_),
    .A3(_0365_),
    .A4(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5138_ (.A1(_0367_),
    .A2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5139_ (.I(_0987_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5140_ (.I(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5141_ (.A1(_0896_),
    .A2(_0982_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5142_ (.A1(_0981_),
    .A2(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5143_ (.A1(_0905_),
    .A2(_0978_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5144_ (.A1(_0905_),
    .A2(_0978_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5145_ (.A1(_0901_),
    .A2(_0992_),
    .A3(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5146_ (.I(_0339_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5147_ (.I(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5148_ (.A1(_0996_),
    .A2(_3299_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5149_ (.A1(_0824_),
    .A2(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5150_ (.A1(_0913_),
    .A2(_0932_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5151_ (.A1(_0909_),
    .A2(_0933_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5152_ (.A1(_0999_),
    .A2(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5153_ (.A1(_0998_),
    .A2(_1001_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5154_ (.I(_0930_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5155_ (.A1(_0923_),
    .A2(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5156_ (.A1(_0917_),
    .A2(_0931_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5157_ (.A1(_1004_),
    .A2(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5158_ (.I(_0946_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5159_ (.A1(_0941_),
    .A2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5160_ (.A1(_0935_),
    .A2(_0936_),
    .B(_0947_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5161_ (.A1(_1008_),
    .A2(_1009_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5162_ (.I(\dspArea_regB[13] ),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5163_ (.I(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5164_ (.I(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5165_ (.A1(_1013_),
    .A2(_0552_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5166_ (.A1(_0332_),
    .A2(_3304_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5167_ (.A1(_0997_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5168_ (.A1(_1014_),
    .A2(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5169_ (.I(\dspArea_regB[10] ),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5170_ (.I(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5171_ (.A1(_1019_),
    .A2(_0670_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5172_ (.A1(_0319_),
    .A2(_0920_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5173_ (.I(_0312_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5174_ (.A1(_1022_),
    .A2(\dspArea_regA[5] ),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5175_ (.A1(_1021_),
    .A2(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5176_ (.A1(_1020_),
    .A2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5177_ (.A1(_0321_),
    .A2(_0433_),
    .A3(_0817_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5178_ (.A1(_0928_),
    .A2(_0466_),
    .A3(_0922_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5179_ (.A1(_1026_),
    .A2(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5180_ (.A1(_1025_),
    .A2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5181_ (.A1(_1017_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5182_ (.A1(_1010_),
    .A2(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5183_ (.A1(_1006_),
    .A2(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5184_ (.I(_0302_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5185_ (.A1(_1033_),
    .A2(_3346_),
    .A3(_0841_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5186_ (.A1(_0942_),
    .A2(_0945_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5187_ (.A1(_1034_),
    .A2(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5188_ (.A1(_0950_),
    .A2(_0952_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5189_ (.I(\dspArea_regA[10] ),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5190_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _5191_ (.A1(_0283_),
    .A2(_0278_),
    .A3(_1039_),
    .A4(_3359_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5192_ (.I(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5193_ (.A1(_0951_),
    .A2(_1037_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5194_ (.A1(_0305_),
    .A2(_0769_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5195_ (.A1(_0300_),
    .A2(_0689_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5196_ (.I(\dspArea_regA[8] ),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5197_ (.A1(_0295_),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5198_ (.A1(_1044_),
    .A2(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5199_ (.A1(_1043_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5200_ (.A1(_1042_),
    .A2(_1048_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5201_ (.A1(_1036_),
    .A2(_1049_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5202_ (.A1(_0624_),
    .A2(_0773_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5203_ (.A1(_0515_),
    .A2(_3366_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5204_ (.A1(_0277_),
    .A2(_0955_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5205_ (.A1(_1052_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5206_ (.A1(_1051_),
    .A2(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5207_ (.I(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5208_ (.A1(_0570_),
    .A2(_3384_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5209_ (.I(\dspArea_regA[13] ),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5210_ (.I(_1058_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5211_ (.A1(_0264_),
    .A2(_1059_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5212_ (.A1(\dspArea_regP[13] ),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5213_ (.A1(_1057_),
    .A2(_1061_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5214_ (.A1(\dspArea_regP[12] ),
    .A2(_0960_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5215_ (.A1(_0957_),
    .A2(_0961_),
    .B(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5216_ (.A1(_1056_),
    .A2(_1062_),
    .A3(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5217_ (.A1(_0962_),
    .A2(_0964_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5218_ (.A1(_0962_),
    .A2(_0964_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5219_ (.A1(_0954_),
    .A2(_1066_),
    .B(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5220_ (.A1(_1065_),
    .A2(_1068_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5221_ (.A1(_1050_),
    .A2(_1069_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5222_ (.A1(_0965_),
    .A2(_0968_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5223_ (.A1(_0948_),
    .A2(_0969_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5224_ (.A1(_1071_),
    .A2(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5225_ (.A1(_1032_),
    .A2(_1070_),
    .A3(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5226_ (.A1(_0971_),
    .A2(_0972_),
    .A3(_0970_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5227_ (.A1(_0971_),
    .A2(_0972_),
    .B(_0970_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5228_ (.A1(_0934_),
    .A2(_1075_),
    .B(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5229_ (.A1(_1074_),
    .A2(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5230_ (.A1(_1002_),
    .A2(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5231_ (.A1(_0974_),
    .A2(_0977_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5232_ (.A1(_1080_),
    .A2(_0993_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5233_ (.A1(_1079_),
    .A2(_1081_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5234_ (.A1(_0994_),
    .A2(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5235_ (.A1(_0991_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5236_ (.I(_0379_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5237_ (.A1(\dspArea_regP[13] ),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5238_ (.I(_0240_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5239_ (.A1(_0989_),
    .A2(_1084_),
    .B(_1086_),
    .C(_1087_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5240_ (.A1(_1079_),
    .A2(_1081_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5241_ (.A1(_0824_),
    .A2(_0997_),
    .A3(_1001_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5242_ (.A1(_1010_),
    .A2(_1030_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5243_ (.A1(_1006_),
    .A2(_1031_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5244_ (.A1(_1090_),
    .A2(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5245_ (.A1(_0995_),
    .A2(_0555_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5246_ (.A1(_0914_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5247_ (.A1(_0350_),
    .A2(_0390_),
    .A3(_1016_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5248_ (.A1(_1094_),
    .A2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5249_ (.A1(_0355_),
    .A2(_0391_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5250_ (.A1(_1096_),
    .A2(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5251_ (.A1(_1092_),
    .A2(_1098_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5252_ (.I(_1028_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5253_ (.A1(_1025_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5254_ (.A1(_1017_),
    .A2(_1029_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5255_ (.A1(_1101_),
    .A2(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5256_ (.I(_1048_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5257_ (.A1(_1042_),
    .A2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5258_ (.A1(_1036_),
    .A2(_1049_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5259_ (.A1(_1105_),
    .A2(_1106_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5260_ (.A1(_0347_),
    .A2(_0461_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5261_ (.I(_0330_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5262_ (.I(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5263_ (.A1(_1110_),
    .A2(_3313_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5264_ (.A1(_1093_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5265_ (.A1(_1108_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5266_ (.A1(_1018_),
    .A2(_3321_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5267_ (.A1(_0735_),
    .A2(\dspArea_regA[5] ),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5268_ (.I(\dspArea_regB[8] ),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5269_ (.A1(_1116_),
    .A2(\dspArea_regA[6] ),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5270_ (.A1(_1115_),
    .A2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5271_ (.A1(_1114_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5272_ (.A1(_0737_),
    .A2(_3330_),
    .A3(_0921_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5273_ (.A1(_1019_),
    .A2(_0670_),
    .A3(_1024_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5274_ (.A1(_1120_),
    .A2(_1121_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5275_ (.A1(_1119_),
    .A2(_1122_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5276_ (.A1(_1113_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5277_ (.A1(_1107_),
    .A2(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5278_ (.A1(_1103_),
    .A2(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5279_ (.A1(_1033_),
    .A2(_3354_),
    .A3(_0944_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5280_ (.A1(_1043_),
    .A2(_1047_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5281_ (.A1(_1127_),
    .A2(_1128_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5282_ (.A1(_0547_),
    .A2(_0956_),
    .A3(_0952_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5283_ (.A1(_0291_),
    .A2(_3360_),
    .A3(_1054_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5284_ (.A1(_0306_),
    .A2(_3345_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5285_ (.A1(_0507_),
    .A2(_1045_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5286_ (.I(\dspArea_regB[5] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5287_ (.A1(_1134_),
    .A2(_3358_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5288_ (.A1(_1133_),
    .A2(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5289_ (.A1(_1132_),
    .A2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5290_ (.A1(_1130_),
    .A2(_1131_),
    .A3(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5291_ (.A1(_1130_),
    .A2(_1131_),
    .B(_1137_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5292_ (.A1(_1138_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5293_ (.A1(_1129_),
    .A2(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5294_ (.A1(_0623_),
    .A2(_1039_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5295_ (.A1(_0514_),
    .A2(_3374_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5296_ (.I(\dspArea_regB[2] ),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5297_ (.A1(_1144_),
    .A2(_0958_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5298_ (.A1(_1143_),
    .A2(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5299_ (.A1(_1142_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5300_ (.I(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5301_ (.I(\dspArea_regB[1] ),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5302_ (.I(_1149_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5303_ (.A1(_1150_),
    .A2(_3390_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5304_ (.A1(_0476_),
    .A2(_3395_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5305_ (.A1(\dspArea_regP[14] ),
    .A2(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5306_ (.A1(_1151_),
    .A2(_1153_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5307_ (.A1(\dspArea_regP[13] ),
    .A2(_1060_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5308_ (.A1(_1057_),
    .A2(_1061_),
    .B(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5309_ (.A1(_1148_),
    .A2(_1154_),
    .A3(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5310_ (.A1(_1062_),
    .A2(_1064_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5311_ (.A1(_1062_),
    .A2(_1064_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5312_ (.A1(_1056_),
    .A2(_1158_),
    .B(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5313_ (.A1(_1157_),
    .A2(_1160_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5314_ (.A1(_1141_),
    .A2(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5315_ (.A1(_1065_),
    .A2(_1068_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5316_ (.A1(_1050_),
    .A2(_1069_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5317_ (.A1(_1163_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5318_ (.A1(_1126_),
    .A2(_1162_),
    .A3(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5319_ (.A1(_1071_),
    .A2(_1072_),
    .A3(_1070_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5320_ (.A1(_1071_),
    .A2(_1072_),
    .B(_1070_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5321_ (.A1(_1032_),
    .A2(_1167_),
    .B(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5322_ (.A1(_1099_),
    .A2(_1166_),
    .A3(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5323_ (.A1(_1074_),
    .A2(_1077_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5324_ (.A1(_1002_),
    .A2(_1078_),
    .B(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5325_ (.A1(_1089_),
    .A2(_1170_),
    .A3(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5326_ (.A1(_1088_),
    .A2(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5327_ (.A1(_0982_),
    .A2(_1083_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5328_ (.A1(_0994_),
    .A2(_0981_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5329_ (.A1(_1082_),
    .A2(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5330_ (.A1(_0897_),
    .A2(_1175_),
    .B(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5331_ (.A1(_1174_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5332_ (.A1(\dspArea_regP[14] ),
    .A2(_0495_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5333_ (.A1(_0451_),
    .A2(_1179_),
    .B(_1180_),
    .C(_1087_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5334_ (.A1(\dspArea_regP[15] ),
    .A2(_0799_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5335_ (.A1(_1170_),
    .A2(_1172_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5336_ (.A1(_1170_),
    .A2(_1172_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5337_ (.A1(_1089_),
    .A2(_1182_),
    .B(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5338_ (.A1(_1092_),
    .A2(_1098_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5339_ (.A1(_1096_),
    .A2(_1097_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5340_ (.A1(_1107_),
    .A2(_1124_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5341_ (.A1(_1103_),
    .A2(_1125_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5342_ (.A1(_1187_),
    .A2(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5343_ (.I(_0342_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5344_ (.A1(_1190_),
    .A2(_3316_),
    .A3(_1015_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5345_ (.A1(_0349_),
    .A2(_0501_),
    .A3(_1112_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5346_ (.A1(_0353_),
    .A2(_0501_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5347_ (.A1(_1191_),
    .A2(_1192_),
    .A3(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5348_ (.A1(_1191_),
    .A2(_1192_),
    .B(_1193_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5349_ (.A1(_1194_),
    .A2(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5350_ (.I(\dspArea_regB[15] ),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5351_ (.I(_1197_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5352_ (.A1(_1198_),
    .A2(_0390_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5353_ (.A1(_1196_),
    .A2(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5354_ (.I(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5355_ (.A1(_1186_),
    .A2(_1189_),
    .A3(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5356_ (.A1(_1119_),
    .A2(_1122_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5357_ (.A1(_1113_),
    .A2(_1123_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5358_ (.A1(_1130_),
    .A2(_1131_),
    .A3(_1137_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5359_ (.A1(_1129_),
    .A2(_1205_),
    .B(_1139_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5360_ (.A1(_1011_),
    .A2(_0555_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5361_ (.A1(_0339_),
    .A2(\dspArea_regA[3] ),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5362_ (.A1(_0330_),
    .A2(_0920_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5363_ (.A1(_1208_),
    .A2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5364_ (.A1(_1207_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5365_ (.A1(_0926_),
    .A2(_0478_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5366_ (.A1(_0318_),
    .A2(\dspArea_regA[6] ),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5367_ (.A1(_0312_),
    .A2(\dspArea_regA[7] ),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5368_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5369_ (.A1(_1212_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5370_ (.A1(_0321_),
    .A2(_3337_),
    .A3(_1023_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5371_ (.A1(_0326_),
    .A2(_0433_),
    .A3(_1118_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5372_ (.A1(_1217_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5373_ (.A1(_1211_),
    .A2(_1216_),
    .A3(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5374_ (.A1(_1206_),
    .A2(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5375_ (.A1(_1203_),
    .A2(_1204_),
    .A3(_1221_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5376_ (.A1(_1203_),
    .A2(_1204_),
    .B(_1221_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5377_ (.A1(_1222_),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5378_ (.I(_0302_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5379_ (.A1(_1225_),
    .A2(_3361_),
    .A3(_1046_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5380_ (.A1(_0308_),
    .A2(_3346_),
    .A3(_1136_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5381_ (.A1(_1226_),
    .A2(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5382_ (.I(_3385_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5383_ (.A1(_0675_),
    .A2(_1229_),
    .A3(_1053_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5384_ (.A1(_0460_),
    .A2(_3369_),
    .A3(_1146_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5385_ (.A1(_0307_),
    .A2(_3354_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5386_ (.I(\dspArea_regB[6] ),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5387_ (.I(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5388_ (.A1(_1234_),
    .A2(_0949_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5389_ (.A1(_0554_),
    .A2(_3366_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5390_ (.A1(_1235_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5391_ (.A1(_1232_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5392_ (.A1(_1230_),
    .A2(_1231_),
    .A3(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5393_ (.A1(_1230_),
    .A2(_1231_),
    .B(_1238_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5394_ (.A1(_1239_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5395_ (.A1(_1228_),
    .A2(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5396_ (.A1(_0768_),
    .A2(_3375_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5397_ (.I(\dspArea_regB[3] ),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5398_ (.A1(_1244_),
    .A2(_0958_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5399_ (.A1(_1144_),
    .A2(\dspArea_regA[13] ),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5400_ (.A1(_1245_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5401_ (.A1(_1243_),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5402_ (.I(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5403_ (.A1(_0694_),
    .A2(_3397_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5404_ (.A1(_0697_),
    .A2(_3404_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5405_ (.A1(\dspArea_regP[15] ),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5406_ (.A1(_1250_),
    .A2(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5407_ (.A1(\dspArea_regP[14] ),
    .A2(_1152_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5408_ (.A1(_1151_),
    .A2(_1153_),
    .B(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5409_ (.A1(_1249_),
    .A2(_1253_),
    .A3(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5410_ (.A1(_1154_),
    .A2(_1156_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5411_ (.A1(_1154_),
    .A2(_1156_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5412_ (.A1(_1148_),
    .A2(_1257_),
    .B(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5413_ (.A1(_1256_),
    .A2(_1259_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5414_ (.A1(_1242_),
    .A2(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5415_ (.A1(_1157_),
    .A2(_1160_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5416_ (.A1(_1141_),
    .A2(_1161_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5417_ (.A1(_1262_),
    .A2(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5418_ (.A1(_1224_),
    .A2(_1261_),
    .A3(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5419_ (.A1(_1163_),
    .A2(_1164_),
    .A3(_1162_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5420_ (.A1(_1163_),
    .A2(_1164_),
    .B(_1162_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5421_ (.A1(_1126_),
    .A2(_1266_),
    .B(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5422_ (.A1(_1202_),
    .A2(_1265_),
    .A3(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5423_ (.A1(_1166_),
    .A2(_1169_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5424_ (.A1(_1166_),
    .A2(_1169_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5425_ (.A1(_1099_),
    .A2(_1270_),
    .B(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5426_ (.A1(_1185_),
    .A2(_1269_),
    .A3(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5427_ (.A1(_1184_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5428_ (.A1(_1088_),
    .A2(_1173_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5429_ (.I(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5430_ (.A1(_1174_),
    .A2(_1178_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5431_ (.A1(_1276_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5432_ (.A1(_1274_),
    .A2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5433_ (.A1(_0989_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5434_ (.A1(_3681_),
    .A2(_1181_),
    .A3(_1280_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5435_ (.I(_1273_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5436_ (.A1(_1184_),
    .A2(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5437_ (.A1(_1174_),
    .A2(_1274_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5438_ (.A1(_1082_),
    .A2(_1176_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5439_ (.A1(_1184_),
    .A2(_1281_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5440_ (.I(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5441_ (.A1(_1275_),
    .A2(_1282_),
    .B1(_1283_),
    .B2(_1284_),
    .C(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5442_ (.A1(_0723_),
    .A2(_0728_),
    .B(_0796_),
    .C(_0878_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5443_ (.A1(_0893_),
    .A2(_0894_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5444_ (.A1(_0982_),
    .A2(_1083_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5445_ (.A1(_1288_),
    .A2(_1289_),
    .B(_1290_),
    .C(_1283_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5446_ (.A1(_1287_),
    .A2(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5447_ (.A1(_1189_),
    .A2(_1201_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5448_ (.A1(_1189_),
    .A2(_1201_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5449_ (.A1(_1186_),
    .A2(_1294_),
    .A3(_1293_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5450_ (.A1(_1293_),
    .A2(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5451_ (.I(_0358_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5452_ (.A1(_1297_),
    .A2(_0391_),
    .A3(_1196_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5453_ (.A1(_1195_),
    .A2(_1298_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5454_ (.I(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5455_ (.A1(_1129_),
    .A2(_1140_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5456_ (.A1(_1139_),
    .A2(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5457_ (.A1(_1302_),
    .A2(_1220_),
    .B(_1223_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5458_ (.A1(_0342_),
    .A2(_3324_),
    .A3(_1111_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5459_ (.I(_1013_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5460_ (.A1(_1305_),
    .A2(_3306_),
    .A3(_1210_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5461_ (.A1(_0352_),
    .A2(_3306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5462_ (.A1(_1304_),
    .A2(_1306_),
    .A3(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5463_ (.A1(_1304_),
    .A2(_1306_),
    .B(_1307_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5464_ (.A1(_1308_),
    .A2(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5465_ (.A1(_1197_),
    .A2(_3301_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5466_ (.A1(_1310_),
    .A2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5467_ (.A1(_1303_),
    .A2(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5468_ (.A1(_1300_),
    .A2(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5469_ (.I(_1219_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5470_ (.A1(_1216_),
    .A2(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5471_ (.A1(_1216_),
    .A2(_1219_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5472_ (.A1(_1211_),
    .A2(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5473_ (.A1(_1230_),
    .A2(_1231_),
    .A3(_1238_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5474_ (.A1(_1228_),
    .A2(_1319_),
    .B(_1240_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5475_ (.A1(_0346_),
    .A2(_0670_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5476_ (.A1(_0340_),
    .A2(_0920_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5477_ (.I(\dspArea_regB[11] ),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5478_ (.A1(_1323_),
    .A2(_3328_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5479_ (.A1(_1322_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5480_ (.A1(_1321_),
    .A2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5481_ (.A1(_0927_),
    .A2(_0769_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5482_ (.A1(_0319_),
    .A2(_0689_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5483_ (.A1(_1022_),
    .A2(_1045_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5484_ (.A1(_1328_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5485_ (.A1(_1327_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5486_ (.A1(_0322_),
    .A2(_0631_),
    .A3(_1117_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5487_ (.I(_0747_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5488_ (.A1(_1333_),
    .A2(_0521_),
    .A3(_1215_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5489_ (.A1(_1332_),
    .A2(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5490_ (.A1(_1326_),
    .A2(_1331_),
    .A3(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5491_ (.A1(_1320_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5492_ (.A1(_1316_),
    .A2(_1318_),
    .A3(_1337_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5493_ (.A1(_1316_),
    .A2(_1318_),
    .B(_1337_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5494_ (.A1(_1338_),
    .A2(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5495_ (.A1(_1033_),
    .A2(_3369_),
    .A3(_1135_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5496_ (.I(_0615_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5497_ (.A1(_1342_),
    .A2(_3354_),
    .A3(_1237_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5498_ (.A1(_1341_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5499_ (.I(_0284_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5500_ (.I(_3390_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5501_ (.A1(_1345_),
    .A2(_1346_),
    .A3(_1145_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5502_ (.I(_0677_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5503_ (.A1(_1348_),
    .A2(_3377_),
    .A3(_1247_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5504_ (.A1(_0551_),
    .A2(_0773_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5505_ (.A1(_0839_),
    .A2(_1039_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5506_ (.I(_0295_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5507_ (.A1(_1352_),
    .A2(_0955_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5508_ (.A1(_1351_),
    .A2(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5509_ (.A1(_1350_),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5510_ (.A1(_1347_),
    .A2(_1349_),
    .A3(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5511_ (.A1(_1347_),
    .A2(_1349_),
    .B(_1355_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5512_ (.A1(_1356_),
    .A2(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5513_ (.A1(_1344_),
    .A2(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5514_ (.A1(_0289_),
    .A2(_0959_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5515_ (.A1(_1244_),
    .A2(_3389_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5516_ (.A1(_0276_),
    .A2(\dspArea_regA[14] ),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5517_ (.A1(_1361_),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5518_ (.A1(_1360_),
    .A2(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5519_ (.I(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5520_ (.A1(_0271_),
    .A2(_3406_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5521_ (.I(\dspArea_regB[0] ),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5522_ (.I(\dspArea_regA[16] ),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5523_ (.A1(_1367_),
    .A2(_1368_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5524_ (.A1(\dspArea_regP[16] ),
    .A2(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5525_ (.A1(_1366_),
    .A2(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5526_ (.A1(\dspArea_regP[15] ),
    .A2(_1251_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5527_ (.A1(_1250_),
    .A2(_1252_),
    .B(_1372_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5528_ (.A1(_1365_),
    .A2(_1371_),
    .A3(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5529_ (.A1(_1253_),
    .A2(_1255_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5530_ (.A1(_1253_),
    .A2(_1255_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5531_ (.A1(_1249_),
    .A2(_1375_),
    .B(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5532_ (.A1(_1374_),
    .A2(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5533_ (.A1(_1359_),
    .A2(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5534_ (.A1(_1256_),
    .A2(_1259_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5535_ (.A1(_1242_),
    .A2(_1260_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5536_ (.A1(_1380_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5537_ (.A1(_1340_),
    .A2(_1379_),
    .A3(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5538_ (.A1(_1262_),
    .A2(_1263_),
    .A3(_1261_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5539_ (.A1(_1262_),
    .A2(_1263_),
    .B(_1261_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5540_ (.A1(_1224_),
    .A2(_1384_),
    .B(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5541_ (.A1(_1314_),
    .A2(_1383_),
    .A3(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5542_ (.A1(_1265_),
    .A2(_1268_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5543_ (.A1(_1265_),
    .A2(_1268_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5544_ (.A1(_1202_),
    .A2(_1388_),
    .B(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5545_ (.A1(_1387_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5546_ (.A1(_1296_),
    .A2(_1391_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5547_ (.A1(_1269_),
    .A2(_1272_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5548_ (.A1(_1269_),
    .A2(_1272_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5549_ (.A1(_1092_),
    .A2(_1098_),
    .A3(_1393_),
    .B(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5550_ (.A1(_1392_),
    .A2(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5551_ (.A1(_1292_),
    .A2(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5552_ (.I0(\dspArea_regP[16] ),
    .I1(_1397_),
    .S(_0726_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5553_ (.A1(_0882_),
    .A2(_1398_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5554_ (.A1(\dspArea_regP[17] ),
    .A2(_0799_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5555_ (.A1(_1387_),
    .A2(_1390_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5556_ (.A1(_1296_),
    .A2(_1391_),
    .B(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5557_ (.A1(_1303_),
    .A2(_1312_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5558_ (.A1(_1300_),
    .A2(_1313_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5559_ (.A1(_1402_),
    .A2(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5560_ (.I(_1297_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5561_ (.I(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5562_ (.I(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5563_ (.A1(_1407_),
    .A2(_3302_),
    .A3(_1310_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5564_ (.A1(_1309_),
    .A2(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5565_ (.A1(_1228_),
    .A2(_1241_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5566_ (.A1(_1240_),
    .A2(_1410_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5567_ (.A1(_1411_),
    .A2(_1336_),
    .B(_1339_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5568_ (.I(_0915_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5569_ (.I(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5570_ (.A1(_1414_),
    .A2(_3332_),
    .A3(_1209_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5571_ (.I(_1305_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5572_ (.A1(_1416_),
    .A2(_3316_),
    .A3(_1325_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5573_ (.I(\dspArea_regB[14] ),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5574_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5575_ (.A1(_1419_),
    .A2(_3316_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5576_ (.A1(_1415_),
    .A2(_1417_),
    .A3(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5577_ (.A1(_1415_),
    .A2(_1417_),
    .B(_1420_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5578_ (.A1(_1421_),
    .A2(_1422_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5579_ (.I(_0358_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5580_ (.A1(_1424_),
    .A2(_3308_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5581_ (.A1(_1423_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5582_ (.A1(_1412_),
    .A2(_1426_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5583_ (.A1(_1409_),
    .A2(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5584_ (.I(_1335_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5585_ (.A1(_1331_),
    .A2(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5586_ (.A1(_1331_),
    .A2(_1335_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5587_ (.A1(_1326_),
    .A2(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5588_ (.A1(_1347_),
    .A2(_1349_),
    .A3(_1355_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5589_ (.A1(_1344_),
    .A2(_1433_),
    .B(_1357_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5590_ (.I(\dspArea_regB[13] ),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5591_ (.A1(_1435_),
    .A2(_3322_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5592_ (.I(\dspArea_regB[12] ),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5593_ (.A1(_1437_),
    .A2(_3328_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5594_ (.A1(_1109_),
    .A2(\dspArea_regA[6] ),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5595_ (.A1(_1438_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5596_ (.A1(_1436_),
    .A2(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5597_ (.A1(_0325_),
    .A2(_3344_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5598_ (.I(\dspArea_regB[9] ),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5599_ (.A1(_1443_),
    .A2(_1045_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5600_ (.I(\dspArea_regB[8] ),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5601_ (.A1(_1445_),
    .A2(\dspArea_regA[9] ),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5602_ (.A1(_1444_),
    .A2(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5603_ (.A1(_1442_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5604_ (.A1(_0924_),
    .A2(_0834_),
    .A3(_1214_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5605_ (.I(_0926_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5606_ (.A1(_1450_),
    .A2(_3337_),
    .A3(_1330_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5607_ (.A1(_1449_),
    .A2(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5608_ (.A1(_1441_),
    .A2(_1448_),
    .A3(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5609_ (.A1(_1434_),
    .A2(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5610_ (.A1(_1430_),
    .A2(_1432_),
    .A3(_1454_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5611_ (.A1(_1430_),
    .A2(_1432_),
    .B(_1454_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5612_ (.A1(_1455_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5613_ (.A1(_0829_),
    .A2(_3377_),
    .A3(_1236_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5614_ (.A1(_0308_),
    .A2(_3361_),
    .A3(_1354_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5615_ (.A1(_1458_),
    .A2(_1459_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5616_ (.A1(_0675_),
    .A2(_3399_),
    .A3(_1246_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5617_ (.A1(_0678_),
    .A2(_1229_),
    .A3(_1363_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5618_ (.A1(_0615_),
    .A2(_3368_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5619_ (.A1(_1234_),
    .A2(_3375_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5620_ (.A1(_0554_),
    .A2(_3383_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5621_ (.A1(_1464_),
    .A2(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5622_ (.A1(_1463_),
    .A2(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5623_ (.A1(_1461_),
    .A2(_1462_),
    .A3(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5624_ (.A1(_1461_),
    .A2(_1462_),
    .B(_1467_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5625_ (.A1(_1468_),
    .A2(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5626_ (.A1(_1460_),
    .A2(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5627_ (.A1(_0768_),
    .A2(_1059_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5628_ (.A1(_1244_),
    .A2(_3395_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5629_ (.A1(_0276_),
    .A2(_3403_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5630_ (.A1(_1473_),
    .A2(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5631_ (.A1(_1472_),
    .A2(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5632_ (.I(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5633_ (.I(_3414_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5634_ (.A1(_0694_),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5635_ (.A1(_0697_),
    .A2(_3422_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5636_ (.A1(\dspArea_regP[17] ),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5637_ (.A1(_1479_),
    .A2(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5638_ (.A1(\dspArea_regP[16] ),
    .A2(_1369_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5639_ (.A1(_1366_),
    .A2(_1370_),
    .B(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5640_ (.A1(_1477_),
    .A2(_1482_),
    .A3(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5641_ (.A1(_1371_),
    .A2(_1373_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5642_ (.A1(_1371_),
    .A2(_1373_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5643_ (.A1(_1365_),
    .A2(_1486_),
    .B(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5644_ (.A1(_1485_),
    .A2(_1488_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5645_ (.A1(_1471_),
    .A2(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5646_ (.A1(_1374_),
    .A2(_1377_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5647_ (.A1(_1359_),
    .A2(_1378_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5648_ (.A1(_1491_),
    .A2(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5649_ (.A1(_1457_),
    .A2(_1490_),
    .A3(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5650_ (.A1(_1380_),
    .A2(_1381_),
    .A3(_1379_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5651_ (.A1(_1380_),
    .A2(_1381_),
    .B(_1379_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5652_ (.A1(_1340_),
    .A2(_1495_),
    .B(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5653_ (.A1(_1494_),
    .A2(_1497_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5654_ (.A1(_1428_),
    .A2(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5655_ (.A1(_1383_),
    .A2(_1386_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5656_ (.A1(_1383_),
    .A2(_1386_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5657_ (.A1(_1314_),
    .A2(_1500_),
    .B(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5658_ (.A1(_1404_),
    .A2(_1499_),
    .A3(_1502_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5659_ (.A1(_1401_),
    .A2(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5660_ (.A1(_1392_),
    .A2(_1395_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5661_ (.I(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5662_ (.I(_1282_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5663_ (.A1(_1174_),
    .A2(_1274_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5664_ (.A1(_1276_),
    .A2(_1507_),
    .B1(_1508_),
    .B2(_1177_),
    .C(_1285_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5665_ (.A1(_0892_),
    .A2(_0895_),
    .B(_1175_),
    .C(_1508_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5666_ (.A1(_1509_),
    .A2(_1510_),
    .B(_1396_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5667_ (.A1(_1506_),
    .A2(_1511_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5668_ (.A1(_1504_),
    .A2(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5669_ (.A1(_0989_),
    .A2(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5670_ (.A1(_3498_),
    .A2(_1399_),
    .A3(_1514_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5671_ (.A1(_1412_),
    .A2(_1426_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5672_ (.I(_1409_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5673_ (.A1(_1516_),
    .A2(_1427_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5674_ (.A1(_1515_),
    .A2(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5675_ (.I(_0359_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5676_ (.A1(_1519_),
    .A2(_3308_),
    .A3(_1423_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5677_ (.A1(_1422_),
    .A2(_1520_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5678_ (.I(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5679_ (.A1(_1344_),
    .A2(_1358_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5680_ (.A1(_1357_),
    .A2(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5681_ (.A1(_1524_),
    .A2(_1453_),
    .B(_1456_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5682_ (.A1(_1413_),
    .A2(_3338_),
    .A3(_1324_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5683_ (.I(_1013_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5684_ (.A1(_1527_),
    .A2(_3325_),
    .A3(_1440_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5685_ (.A1(_1418_),
    .A2(_3325_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5686_ (.A1(_1526_),
    .A2(_1528_),
    .A3(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5687_ (.A1(_1526_),
    .A2(_1528_),
    .B(_1529_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5688_ (.A1(_1530_),
    .A2(_1531_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5689_ (.I(_1197_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5690_ (.A1(_1533_),
    .A2(_3317_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5691_ (.A1(_1532_),
    .A2(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5692_ (.A1(_1525_),
    .A2(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5693_ (.A1(_1522_),
    .A2(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5694_ (.I(_1452_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5695_ (.A1(_1448_),
    .A2(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5696_ (.A1(_1448_),
    .A2(_1452_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5697_ (.A1(_1441_),
    .A2(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5698_ (.A1(_1461_),
    .A2(_1462_),
    .A3(_1467_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5699_ (.A1(_1460_),
    .A2(_1542_),
    .B(_1469_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5700_ (.A1(_0346_),
    .A2(_3330_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5701_ (.A1(_0340_),
    .A2(_3335_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5702_ (.A1(_0331_),
    .A2(_3343_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5703_ (.A1(_1545_),
    .A2(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5704_ (.A1(_1544_),
    .A2(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5705_ (.A1(_1019_),
    .A2(_0695_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5706_ (.A1(_0319_),
    .A2(_3358_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5707_ (.A1(_1022_),
    .A2(_1038_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5708_ (.A1(_1550_),
    .A2(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5709_ (.A1(_1549_),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5710_ (.A1(_0322_),
    .A2(_3360_),
    .A3(_1329_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5711_ (.A1(_1333_),
    .A2(_3346_),
    .A3(_1447_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5712_ (.A1(_1554_),
    .A2(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5713_ (.A1(_1548_),
    .A2(_1553_),
    .A3(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5714_ (.A1(_1543_),
    .A2(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5715_ (.A1(_1539_),
    .A2(_1541_),
    .A3(_1558_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5716_ (.A1(_1539_),
    .A2(_1541_),
    .B(_1558_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5717_ (.A1(_1559_),
    .A2(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5718_ (.A1(_1033_),
    .A2(_1229_),
    .A3(_1353_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5719_ (.A1(_1342_),
    .A2(_3369_),
    .A3(_1466_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5720_ (.A1(_1562_),
    .A2(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5721_ (.A1(_1345_),
    .A2(_3408_),
    .A3(_1362_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5722_ (.A1(_1348_),
    .A2(_1346_),
    .A3(_1475_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5723_ (.A1(_0551_),
    .A2(_3376_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5724_ (.A1(_0507_),
    .A2(_0959_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5725_ (.A1(_0296_),
    .A2(_1059_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5726_ (.A1(_1568_),
    .A2(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5727_ (.A1(_1567_),
    .A2(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5728_ (.A1(_1565_),
    .A2(_1566_),
    .A3(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5729_ (.A1(_1565_),
    .A2(_1566_),
    .B(_1571_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5730_ (.A1(_1572_),
    .A2(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5731_ (.A1(_1564_),
    .A2(_1574_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5732_ (.A1(_0623_),
    .A2(_3396_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5733_ (.A1(_0514_),
    .A2(_3404_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5734_ (.A1(_1144_),
    .A2(_1368_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5735_ (.A1(_1577_),
    .A2(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5736_ (.A1(_1576_),
    .A2(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5737_ (.I(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5738_ (.I(_3422_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5739_ (.A1(_1150_),
    .A2(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5740_ (.A1(_0476_),
    .A2(\dspArea_regA[18] ),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5741_ (.A1(\dspArea_regP[18] ),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5742_ (.A1(_1583_),
    .A2(_1585_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5743_ (.A1(\dspArea_regP[17] ),
    .A2(_1480_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5744_ (.A1(_1479_),
    .A2(_1481_),
    .B(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5745_ (.A1(_1581_),
    .A2(_1586_),
    .A3(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5746_ (.A1(_1482_),
    .A2(_1484_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5747_ (.A1(_1482_),
    .A2(_1484_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5748_ (.A1(_1477_),
    .A2(_1590_),
    .B(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5749_ (.A1(_1589_),
    .A2(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5750_ (.A1(_1575_),
    .A2(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5751_ (.A1(_1485_),
    .A2(_1488_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5752_ (.A1(_1471_),
    .A2(_1489_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5753_ (.A1(_1595_),
    .A2(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5754_ (.A1(_1561_),
    .A2(_1594_),
    .A3(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5755_ (.A1(_1491_),
    .A2(_1492_),
    .A3(_1490_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5756_ (.A1(_1491_),
    .A2(_1492_),
    .B(_1490_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5757_ (.A1(_1457_),
    .A2(_1599_),
    .B(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5758_ (.A1(_1537_),
    .A2(_1598_),
    .A3(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5759_ (.A1(_1494_),
    .A2(_1497_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5760_ (.A1(_1428_),
    .A2(_1498_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5761_ (.A1(_1603_),
    .A2(_1604_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5762_ (.A1(_1518_),
    .A2(_1602_),
    .A3(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5763_ (.A1(_1499_),
    .A2(_1502_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5764_ (.A1(_1499_),
    .A2(_1502_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5765_ (.A1(_1404_),
    .A2(_1607_),
    .B(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5766_ (.A1(_1606_),
    .A2(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5767_ (.A1(_1396_),
    .A2(_1504_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5768_ (.A1(_1296_),
    .A2(_1391_),
    .B(_1503_),
    .C(_1400_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5769_ (.A1(_1392_),
    .A2(_1395_),
    .A3(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5770_ (.A1(_1404_),
    .A2(_1607_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5771_ (.A1(_1404_),
    .A2(_1607_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5772_ (.A1(_1401_),
    .A2(_1614_),
    .A3(_1615_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5773_ (.A1(_1292_),
    .A2(_1611_),
    .B(_1613_),
    .C(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5774_ (.A1(_1610_),
    .A2(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5775_ (.I(_0395_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5776_ (.I0(\dspArea_regP[18] ),
    .I1(_1618_),
    .S(_1619_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5777_ (.A1(_0882_),
    .A2(_1620_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5778_ (.A1(_1603_),
    .A2(_1604_),
    .A3(_1602_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5779_ (.A1(_1603_),
    .A2(_1604_),
    .B(_1602_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5780_ (.A1(_1518_),
    .A2(_1621_),
    .B(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5781_ (.A1(_1525_),
    .A2(_1535_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5782_ (.A1(_1522_),
    .A2(_1536_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5783_ (.A1(_1624_),
    .A2(_1625_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5784_ (.A1(_1406_),
    .A2(_3317_),
    .A3(_1532_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5785_ (.A1(_1531_),
    .A2(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5786_ (.A1(_1460_),
    .A2(_1470_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5787_ (.A1(_1469_),
    .A2(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5788_ (.A1(_1630_),
    .A2(_1557_),
    .B(_1560_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5789_ (.I(_0915_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5790_ (.A1(_1632_),
    .A2(_3347_),
    .A3(_1439_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5791_ (.I(_0348_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5792_ (.A1(_1634_),
    .A2(_3332_),
    .A3(_1547_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5793_ (.I(_0352_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5794_ (.A1(_1636_),
    .A2(_3332_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5795_ (.A1(_1633_),
    .A2(_1635_),
    .A3(_1637_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5796_ (.A1(_1633_),
    .A2(_1635_),
    .B(_1637_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5797_ (.A1(_1638_),
    .A2(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5798_ (.A1(_1198_),
    .A2(_3326_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5799_ (.A1(_1640_),
    .A2(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5800_ (.A1(_1631_),
    .A2(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5801_ (.A1(_1628_),
    .A2(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5802_ (.I(_1556_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5803_ (.A1(_1553_),
    .A2(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5804_ (.A1(_1553_),
    .A2(_1556_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5805_ (.A1(_1548_),
    .A2(_1647_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5806_ (.A1(_1565_),
    .A2(_1566_),
    .A3(_1571_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5807_ (.A1(_1564_),
    .A2(_1649_),
    .B(_1573_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5808_ (.A1(_1435_),
    .A2(_0769_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5809_ (.A1(_0339_),
    .A2(_3343_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5810_ (.A1(_1109_),
    .A2(\dspArea_regA[8] ),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5811_ (.A1(_1652_),
    .A2(_1653_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5812_ (.A1(_1651_),
    .A2(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5813_ (.A1(_0325_),
    .A2(_0949_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5814_ (.A1(_0735_),
    .A2(\dspArea_regA[10] ),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5815_ (.A1(_1116_),
    .A2(\dspArea_regA[11] ),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5816_ (.A1(_1657_),
    .A2(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5817_ (.A1(_1656_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5818_ (.A1(_0924_),
    .A2(_3367_),
    .A3(_1446_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5819_ (.A1(_1450_),
    .A2(_0834_),
    .A3(_1552_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5820_ (.A1(_1661_),
    .A2(_1662_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5821_ (.A1(_1655_),
    .A2(_1660_),
    .A3(_1663_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5822_ (.A1(_1650_),
    .A2(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5823_ (.A1(_1646_),
    .A2(_1648_),
    .A3(_1665_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5824_ (.A1(_1646_),
    .A2(_1648_),
    .B(_1665_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5825_ (.A1(_1666_),
    .A2(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5826_ (.A1(_0302_),
    .A2(_3391_),
    .A3(_1465_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5827_ (.A1(_0307_),
    .A2(_0956_),
    .A3(_1570_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5828_ (.A1(_1669_),
    .A2(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5829_ (.A1(_0465_),
    .A2(_1478_),
    .A3(_1474_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5830_ (.A1(_0290_),
    .A2(_3397_),
    .A3(_1579_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5831_ (.A1(\dspArea_regB[7] ),
    .A2(_0959_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5832_ (.A1(\dspArea_regB[6] ),
    .A2(_3389_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5833_ (.I(\dspArea_regA[14] ),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5834_ (.A1(_0295_),
    .A2(_1676_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5835_ (.A1(_1675_),
    .A2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5836_ (.A1(_1674_),
    .A2(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5837_ (.A1(_1672_),
    .A2(_1673_),
    .A3(_1679_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5838_ (.A1(_1672_),
    .A2(_1673_),
    .B(_1679_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5839_ (.A1(_1680_),
    .A2(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5840_ (.A1(_1671_),
    .A2(_1682_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5841_ (.A1(_0622_),
    .A2(_3405_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5842_ (.A1(\dspArea_regB[3] ),
    .A2(_1368_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5843_ (.A1(\dspArea_regB[2] ),
    .A2(\dspArea_regA[17] ),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5844_ (.A1(_1685_),
    .A2(_1686_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5845_ (.A1(_1684_),
    .A2(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5846_ (.I(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5847_ (.A1(_0271_),
    .A2(_3432_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5848_ (.A1(_1367_),
    .A2(\dspArea_regA[19] ),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5849_ (.A1(\dspArea_regP[19] ),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5850_ (.A1(_1690_),
    .A2(_1692_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5851_ (.A1(\dspArea_regP[18] ),
    .A2(_1584_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5852_ (.A1(_1583_),
    .A2(_1585_),
    .B(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5853_ (.A1(_1689_),
    .A2(_1693_),
    .A3(_1695_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5854_ (.A1(_1586_),
    .A2(_1588_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5855_ (.A1(_1586_),
    .A2(_1588_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5856_ (.A1(_1581_),
    .A2(_1697_),
    .B(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5857_ (.A1(_1683_),
    .A2(_1696_),
    .A3(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5858_ (.A1(_1589_),
    .A2(_1592_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5859_ (.A1(_1575_),
    .A2(_1593_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5860_ (.A1(_1701_),
    .A2(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5861_ (.A1(_1668_),
    .A2(_1700_),
    .A3(_1703_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5862_ (.A1(_1595_),
    .A2(_1596_),
    .A3(_1594_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5863_ (.A1(_1595_),
    .A2(_1596_),
    .B(_1594_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5864_ (.A1(_1561_),
    .A2(_1705_),
    .B(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5865_ (.A1(_1704_),
    .A2(_1707_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5866_ (.A1(_1644_),
    .A2(_1708_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5867_ (.A1(_1598_),
    .A2(_1601_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5868_ (.A1(_1598_),
    .A2(_1601_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5869_ (.A1(_1537_),
    .A2(_1710_),
    .B(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5870_ (.A1(_1709_),
    .A2(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5871_ (.A1(_1626_),
    .A2(_1713_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5872_ (.A1(_1623_),
    .A2(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5873_ (.A1(_1606_),
    .A2(_1609_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5874_ (.A1(_1606_),
    .A2(_1609_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5875_ (.A1(_1717_),
    .A2(_1617_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5876_ (.A1(_1716_),
    .A2(_1718_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5877_ (.A1(_1715_),
    .A2(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5878_ (.A1(\dspArea_regP[19] ),
    .A2(_1085_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5879_ (.A1(_0989_),
    .A2(_1720_),
    .B(_1721_),
    .C(_1087_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5880_ (.A1(_1631_),
    .A2(_1642_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5881_ (.I(_1628_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5882_ (.A1(_1723_),
    .A2(_1643_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5883_ (.A1(_1722_),
    .A2(_1724_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5884_ (.A1(_1406_),
    .A2(_3326_),
    .A3(_1640_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5885_ (.A1(_1639_),
    .A2(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5886_ (.I(_1727_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5887_ (.A1(_1564_),
    .A2(_1574_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5888_ (.A1(_1573_),
    .A2(_1729_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5889_ (.A1(_1730_),
    .A2(_1664_),
    .B(_1667_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5890_ (.A1(_1190_),
    .A2(_3355_),
    .A3(_1546_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5891_ (.A1(_1416_),
    .A2(_3339_),
    .A3(_1654_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5892_ (.A1(_0353_),
    .A2(_3339_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5893_ (.A1(_1732_),
    .A2(_1733_),
    .A3(_1734_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5894_ (.A1(_1732_),
    .A2(_1733_),
    .B(_1734_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5895_ (.A1(_1735_),
    .A2(_1736_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5896_ (.A1(_1198_),
    .A2(_3333_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5897_ (.A1(_1737_),
    .A2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5898_ (.A1(_1731_),
    .A2(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5899_ (.A1(_1728_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5900_ (.I(_1663_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5901_ (.A1(_1660_),
    .A2(_1742_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5902_ (.A1(_1660_),
    .A2(_1663_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5903_ (.A1(_1655_),
    .A2(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5904_ (.A1(_1672_),
    .A2(_1673_),
    .A3(_1679_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5905_ (.A1(_1671_),
    .A2(_1746_),
    .B(_1681_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5906_ (.A1(_1012_),
    .A2(_0631_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5907_ (.A1(_0995_),
    .A2(_3352_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5908_ (.A1(_1110_),
    .A2(_0949_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5909_ (.A1(_1749_),
    .A2(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5910_ (.A1(_1748_),
    .A2(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5911_ (.A1(_0326_),
    .A2(_3367_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5912_ (.A1(_0736_),
    .A2(_0955_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5913_ (.I(_1116_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5914_ (.A1(_1755_),
    .A2(_3383_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5915_ (.A1(_1754_),
    .A2(_1756_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5916_ (.A1(_1753_),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5917_ (.I(_0737_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5918_ (.A1(_1759_),
    .A2(_3377_),
    .A3(_1551_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5919_ (.A1(_0748_),
    .A2(_3361_),
    .A3(_1659_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5920_ (.A1(_1760_),
    .A2(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5921_ (.A1(_1752_),
    .A2(_1758_),
    .A3(_1762_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5922_ (.A1(_1747_),
    .A2(_1763_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5923_ (.A1(_1743_),
    .A2(_1745_),
    .A3(_1764_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5924_ (.A1(_1743_),
    .A2(_1745_),
    .B(_1764_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5925_ (.A1(_1765_),
    .A2(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5926_ (.A1(_0829_),
    .A2(_3399_),
    .A3(_1569_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5927_ (.A1(_0608_),
    .A2(_1229_),
    .A3(_1678_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5928_ (.A1(_1768_),
    .A2(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5929_ (.A1(_0285_),
    .A2(_3425_),
    .A3(_1578_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5930_ (.A1(_0460_),
    .A2(_3408_),
    .A3(_1687_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5931_ (.A1(_0307_),
    .A2(_3391_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5932_ (.A1(_1234_),
    .A2(_3396_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5933_ (.I(_1134_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5934_ (.A1(_1775_),
    .A2(_3405_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5935_ (.A1(_1774_),
    .A2(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5936_ (.A1(_1773_),
    .A2(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5937_ (.A1(_1771_),
    .A2(_1772_),
    .A3(_1778_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5938_ (.A1(_1771_),
    .A2(_1772_),
    .B(_1778_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5939_ (.A1(_1779_),
    .A2(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5940_ (.A1(_1770_),
    .A2(_1781_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5941_ (.A1(_0562_),
    .A2(_3415_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5942_ (.A1(_0564_),
    .A2(_3423_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5943_ (.A1(_0469_),
    .A2(_3431_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5944_ (.A1(_1784_),
    .A2(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5945_ (.A1(_1783_),
    .A2(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5946_ (.A1(_1149_),
    .A2(_3439_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5947_ (.A1(_0263_),
    .A2(_3447_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5948_ (.A1(\dspArea_regP[20] ),
    .A2(_1789_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5949_ (.A1(_1788_),
    .A2(_1790_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5950_ (.A1(\dspArea_regP[19] ),
    .A2(_1691_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5951_ (.A1(_1690_),
    .A2(_1692_),
    .B(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5952_ (.A1(_1791_),
    .A2(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5953_ (.A1(_1787_),
    .A2(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5954_ (.A1(_1693_),
    .A2(_1695_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5955_ (.A1(_1693_),
    .A2(_1695_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5956_ (.A1(_1689_),
    .A2(_1796_),
    .B(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5957_ (.A1(_1795_),
    .A2(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5958_ (.A1(_1782_),
    .A2(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5959_ (.A1(_1696_),
    .A2(_1699_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5960_ (.A1(_1696_),
    .A2(_1699_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5961_ (.A1(_1683_),
    .A2(_1801_),
    .B(_1802_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5962_ (.A1(_1800_),
    .A2(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5963_ (.A1(_1767_),
    .A2(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5964_ (.A1(_1701_),
    .A2(_1702_),
    .A3(_1700_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5965_ (.A1(_1701_),
    .A2(_1702_),
    .B(_1700_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5966_ (.A1(_1668_),
    .A2(_1806_),
    .B(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5967_ (.A1(_1741_),
    .A2(_1805_),
    .A3(_1808_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5968_ (.A1(_1704_),
    .A2(_1707_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5969_ (.A1(_1644_),
    .A2(_1708_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5970_ (.A1(_1810_),
    .A2(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5971_ (.A1(_1725_),
    .A2(_1809_),
    .A3(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5972_ (.A1(_1709_),
    .A2(_1712_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5973_ (.A1(_1626_),
    .A2(_1713_),
    .B(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5974_ (.A1(_1813_),
    .A2(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5975_ (.A1(_1813_),
    .A2(_1815_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5976_ (.A1(_1816_),
    .A2(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5977_ (.A1(_1623_),
    .A2(_1714_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5978_ (.A1(_1623_),
    .A2(_1714_),
    .B(_1606_),
    .C(_1609_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5979_ (.A1(_1819_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5980_ (.A1(_1616_),
    .A2(_1613_),
    .B(_1715_),
    .C(_1610_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5981_ (.A1(_1623_),
    .A2(_1714_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5982_ (.A1(_1717_),
    .A2(_1823_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5983_ (.I(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5984_ (.A1(_1287_),
    .A2(_1291_),
    .B(_1611_),
    .C(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5985_ (.A1(_1821_),
    .A2(_1822_),
    .A3(_1826_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5986_ (.A1(_1818_),
    .A2(_1827_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5987_ (.I0(\dspArea_regP[20] ),
    .I1(_1828_),
    .S(_1619_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5988_ (.A1(_0882_),
    .A2(_1829_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5989_ (.I(\dspArea_regP[21] ),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5990_ (.I(_0987_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5991_ (.A1(_1818_),
    .A2(_1827_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5992_ (.A1(_1810_),
    .A2(_1811_),
    .A3(_1809_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5993_ (.A1(_1810_),
    .A2(_1811_),
    .B(_1809_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5994_ (.A1(_1725_),
    .A2(_1833_),
    .B(_1834_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5995_ (.A1(_1731_),
    .A2(_1739_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5996_ (.A1(_1728_),
    .A2(_1740_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5997_ (.A1(_1836_),
    .A2(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5998_ (.A1(_1407_),
    .A2(_3333_),
    .A3(_1737_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5999_ (.A1(_1736_),
    .A2(_1839_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6000_ (.A1(_1671_),
    .A2(_1682_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6001_ (.A1(_1681_),
    .A2(_1841_),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6002_ (.A1(_1842_),
    .A2(_1763_),
    .B(_1766_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6003_ (.A1(_1414_),
    .A2(_3362_),
    .A3(_1653_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6004_ (.I(_0348_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6005_ (.A1(_1845_),
    .A2(_3347_),
    .A3(_1751_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6006_ (.I(_1418_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6007_ (.A1(_1847_),
    .A2(_3347_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6008_ (.A1(_1844_),
    .A2(_1846_),
    .A3(_1848_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6009_ (.A1(_1844_),
    .A2(_1846_),
    .B(_1848_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6010_ (.A1(_1849_),
    .A2(_1850_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6011_ (.A1(_0359_),
    .A2(_3340_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6012_ (.A1(_1851_),
    .A2(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6013_ (.A1(_1843_),
    .A2(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6014_ (.A1(_1840_),
    .A2(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6015_ (.I(_1762_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6016_ (.A1(_1758_),
    .A2(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6017_ (.A1(_1758_),
    .A2(_1762_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6018_ (.A1(_1752_),
    .A2(_1858_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6019_ (.A1(_1771_),
    .A2(_1772_),
    .A3(_1778_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6020_ (.A1(_1770_),
    .A2(_1860_),
    .B(_1780_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6021_ (.A1(_1012_),
    .A2(_3353_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6022_ (.A1(_0340_),
    .A2(_3358_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6023_ (.A1(_0331_),
    .A2(_1038_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6024_ (.A1(_1863_),
    .A2(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6025_ (.A1(_1862_),
    .A2(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6026_ (.A1(_1019_),
    .A2(_3376_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6027_ (.A1(_0815_),
    .A2(_0958_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6028_ (.A1(_1022_),
    .A2(_3389_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6029_ (.A1(_1868_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6030_ (.A1(_1867_),
    .A2(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6031_ (.A1(_0322_),
    .A2(_3385_),
    .A3(_1658_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6032_ (.A1(_1333_),
    .A2(_3368_),
    .A3(_1757_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6033_ (.A1(_1872_),
    .A2(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6034_ (.A1(_1866_),
    .A2(_1871_),
    .A3(_1874_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6035_ (.A1(_1861_),
    .A2(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6036_ (.A1(_1857_),
    .A2(_1859_),
    .A3(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6037_ (.A1(_1857_),
    .A2(_1859_),
    .B(_1876_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6038_ (.A1(_1877_),
    .A2(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6039_ (.A1(_1225_),
    .A2(_3408_),
    .A3(_1677_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6040_ (.A1(_0308_),
    .A2(_1346_),
    .A3(_1777_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6041_ (.A1(_1880_),
    .A2(_1881_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6042_ (.A1(_0675_),
    .A2(_3433_),
    .A3(_1686_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6043_ (.I(_1478_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6044_ (.A1(_0678_),
    .A2(_1884_),
    .A3(_1786_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6045_ (.I(_0614_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6046_ (.A1(_1886_),
    .A2(_3398_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6047_ (.A1(_0604_),
    .A2(_3405_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6048_ (.A1(_1352_),
    .A2(_3413_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6049_ (.A1(_1888_),
    .A2(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6050_ (.A1(_1887_),
    .A2(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6051_ (.A1(_1883_),
    .A2(_1885_),
    .A3(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6052_ (.A1(_1883_),
    .A2(_1885_),
    .B(_1891_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6053_ (.A1(_1892_),
    .A2(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6054_ (.A1(_1882_),
    .A2(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6055_ (.A1(_0623_),
    .A2(_1582_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6056_ (.A1(_0514_),
    .A2(_3431_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6057_ (.A1(_1144_),
    .A2(_3438_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6058_ (.A1(_1897_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6059_ (.A1(_1896_),
    .A2(_1899_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6060_ (.A1(_0694_),
    .A2(_3448_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6061_ (.A1(_0697_),
    .A2(\dspArea_regA[21] ),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6062_ (.A1(\dspArea_regP[21] ),
    .A2(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6063_ (.A1(_1901_),
    .A2(_1903_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6064_ (.A1(\dspArea_regP[20] ),
    .A2(_1789_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6065_ (.A1(_1788_),
    .A2(_1790_),
    .B(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6066_ (.A1(_1900_),
    .A2(_1904_),
    .A3(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6067_ (.I(_1787_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6068_ (.A1(_1791_),
    .A2(_1793_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6069_ (.A1(_1791_),
    .A2(_1793_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6070_ (.A1(_1908_),
    .A2(_1909_),
    .B(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6071_ (.A1(_1907_),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6072_ (.A1(_1895_),
    .A2(_1912_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6073_ (.A1(_1787_),
    .A2(_1794_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6074_ (.A1(_1787_),
    .A2(_1794_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6075_ (.A1(_1914_),
    .A2(_1915_),
    .A3(_1798_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6076_ (.A1(_1782_),
    .A2(_1799_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6077_ (.A1(_1916_),
    .A2(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6078_ (.A1(_1879_),
    .A2(_1913_),
    .A3(_1918_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6079_ (.A1(_1800_),
    .A2(_1803_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6080_ (.A1(_1767_),
    .A2(_1804_),
    .B(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6081_ (.A1(_1919_),
    .A2(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6082_ (.A1(_1855_),
    .A2(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6083_ (.A1(_1805_),
    .A2(_1808_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6084_ (.A1(_1805_),
    .A2(_1808_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6085_ (.A1(_1741_),
    .A2(_1924_),
    .B(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6086_ (.A1(_1838_),
    .A2(_1923_),
    .A3(_1926_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6087_ (.A1(_1835_),
    .A2(_1927_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6088_ (.A1(_1817_),
    .A2(_1832_),
    .A3(_1928_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6089_ (.A1(_1817_),
    .A2(_1832_),
    .B(_1928_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6090_ (.A1(_1831_),
    .A2(_1929_),
    .A3(_1930_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6091_ (.A1(_1830_),
    .A2(_0424_),
    .B(_1931_),
    .C(_1087_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6092_ (.I(_3558_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6093_ (.A1(_1843_),
    .A2(_1853_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6094_ (.I(_1840_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6095_ (.A1(_1934_),
    .A2(_1854_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6096_ (.A1(_1933_),
    .A2(_1935_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6097_ (.A1(_1407_),
    .A2(_3340_),
    .A3(_1851_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6098_ (.A1(_1850_),
    .A2(_1937_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6099_ (.A1(_1770_),
    .A2(_1781_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6100_ (.A1(_1780_),
    .A2(_1939_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6101_ (.A1(_1940_),
    .A2(_1875_),
    .B(_1878_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6102_ (.A1(_1190_),
    .A2(_3370_),
    .A3(_1750_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6103_ (.A1(_1416_),
    .A2(_3355_),
    .A3(_1865_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6104_ (.A1(_1419_),
    .A2(_3355_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6105_ (.A1(_1942_),
    .A2(_1943_),
    .A3(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6106_ (.A1(_1942_),
    .A2(_1943_),
    .B(_1944_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6107_ (.A1(_1945_),
    .A2(_1946_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6108_ (.A1(_1424_),
    .A2(_3348_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6109_ (.A1(_1947_),
    .A2(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6110_ (.A1(_1941_),
    .A2(_1949_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6111_ (.A1(_1938_),
    .A2(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6112_ (.I(_1874_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6113_ (.A1(_1871_),
    .A2(_1952_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6114_ (.A1(_1871_),
    .A2(_1874_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6115_ (.A1(_1866_),
    .A2(_1954_),
    .Z(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6116_ (.A1(_1883_),
    .A2(_1885_),
    .A3(_1891_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6117_ (.A1(_1882_),
    .A2(_1956_),
    .B(_1893_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6118_ (.A1(_0346_),
    .A2(_3359_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6119_ (.A1(_1437_),
    .A2(_1038_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6120_ (.A1(_1323_),
    .A2(_3374_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6121_ (.A1(_1959_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6122_ (.A1(_1958_),
    .A2(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6123_ (.A1(_0927_),
    .A2(_3384_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6124_ (.A1(_1443_),
    .A2(_1058_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6125_ (.A1(_1445_),
    .A2(_1676_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6126_ (.A1(_1964_),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6127_ (.A1(_1963_),
    .A2(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6128_ (.I(_0320_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6129_ (.A1(_1968_),
    .A2(_3391_),
    .A3(_1756_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6130_ (.I(_1018_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6131_ (.A1(_1970_),
    .A2(_0956_),
    .A3(_1870_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6132_ (.A1(_1969_),
    .A2(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6133_ (.A1(_1962_),
    .A2(_1967_),
    .A3(_1972_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6134_ (.A1(_1957_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6135_ (.A1(_1953_),
    .A2(_1955_),
    .A3(_1974_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6136_ (.A1(_1953_),
    .A2(_1955_),
    .B(_1974_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6137_ (.A1(_1975_),
    .A2(_1976_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6138_ (.A1(_1225_),
    .A2(_1884_),
    .A3(_1776_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6139_ (.A1(_1342_),
    .A2(_3399_),
    .A3(_1890_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6140_ (.A1(_1978_),
    .A2(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6141_ (.A1(_1345_),
    .A2(_3442_),
    .A3(_1785_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6142_ (.A1(_1348_),
    .A2(_3425_),
    .A3(_1899_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6143_ (.A1(_1886_),
    .A2(_3407_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6144_ (.A1(_0839_),
    .A2(_3414_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6145_ (.A1(_1352_),
    .A2(_3422_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6146_ (.A1(_1984_),
    .A2(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6147_ (.A1(_1983_),
    .A2(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6148_ (.A1(_1981_),
    .A2(_1982_),
    .A3(_1987_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6149_ (.A1(_1981_),
    .A2(_1982_),
    .B(_1987_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6150_ (.A1(_1988_),
    .A2(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6151_ (.A1(_1980_),
    .A2(_1990_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6152_ (.I(_3431_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6153_ (.A1(_0289_),
    .A2(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6154_ (.A1(_1244_),
    .A2(\dspArea_regA[19] ),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6155_ (.A1(_0276_),
    .A2(\dspArea_regA[20] ),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6156_ (.A1(_1994_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6157_ (.A1(_1993_),
    .A2(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6158_ (.I(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6159_ (.A1(_0271_),
    .A2(_3456_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6160_ (.A1(_1367_),
    .A2(\dspArea_regA[22] ),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6161_ (.A1(\dspArea_regP[22] ),
    .A2(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6162_ (.A1(_1999_),
    .A2(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6163_ (.A1(\dspArea_regP[21] ),
    .A2(_1902_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6164_ (.A1(_1901_),
    .A2(_1903_),
    .B(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6165_ (.A1(_1998_),
    .A2(_2002_),
    .A3(_2004_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6166_ (.I(_1900_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6167_ (.A1(_1904_),
    .A2(_1906_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6168_ (.A1(_1904_),
    .A2(_1906_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6169_ (.A1(_2006_),
    .A2(_2007_),
    .B(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6170_ (.A1(_2005_),
    .A2(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6171_ (.A1(_1991_),
    .A2(_2010_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6172_ (.A1(_1910_),
    .A2(_1915_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6173_ (.A1(_1907_),
    .A2(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6174_ (.A1(_1895_),
    .A2(_1912_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6175_ (.A1(_2013_),
    .A2(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6176_ (.A1(_1977_),
    .A2(_2011_),
    .A3(_2015_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6177_ (.A1(_1916_),
    .A2(_1917_),
    .A3(_1913_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6178_ (.A1(_1916_),
    .A2(_1917_),
    .B(_1913_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6179_ (.A1(_1879_),
    .A2(_2017_),
    .B(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6180_ (.A1(_2016_),
    .A2(_2019_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6181_ (.A1(_1951_),
    .A2(_2020_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6182_ (.A1(_1767_),
    .A2(_1804_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6183_ (.A1(_1920_),
    .A2(_2022_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6184_ (.A1(_1919_),
    .A2(_2023_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6185_ (.A1(_1855_),
    .A2(_1922_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6186_ (.A1(_2024_),
    .A2(_2025_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6187_ (.A1(_1936_),
    .A2(_2021_),
    .A3(_2026_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6188_ (.A1(_1923_),
    .A2(_1926_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6189_ (.A1(_1923_),
    .A2(_1926_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6190_ (.A1(_1838_),
    .A2(_2028_),
    .B(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6191_ (.A1(_2027_),
    .A2(_2030_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6192_ (.A1(_1838_),
    .A2(_2028_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6193_ (.A1(_1838_),
    .A2(_2028_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6194_ (.A1(_1835_),
    .A2(_2032_),
    .A3(_2033_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6195_ (.A1(_1725_),
    .A2(_1833_),
    .B(_1834_),
    .C(_1927_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6196_ (.A1(_1813_),
    .A2(_1815_),
    .A3(_2035_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6197_ (.A1(_2034_),
    .A2(_2036_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6198_ (.I(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6199_ (.A1(_1816_),
    .A2(_1817_),
    .A3(_1928_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6200_ (.A1(_1821_),
    .A2(_1822_),
    .A3(_1826_),
    .B(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6201_ (.A1(_2038_),
    .A2(_2040_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6202_ (.A1(_2031_),
    .A2(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6203_ (.I0(\dspArea_regP[22] ),
    .I1(_2042_),
    .S(_1619_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6204_ (.A1(_1932_),
    .A2(_2043_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6205_ (.A1(\dspArea_regP[23] ),
    .A2(_1085_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6206_ (.I(_1831_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6207_ (.A1(_2024_),
    .A2(_2025_),
    .A3(_2021_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6208_ (.A1(_2024_),
    .A2(_2025_),
    .B(_2021_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6209_ (.A1(_1936_),
    .A2(_2046_),
    .B(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6210_ (.A1(_1941_),
    .A2(_1949_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6211_ (.I(_1938_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6212_ (.A1(_2050_),
    .A2(_1950_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6213_ (.A1(_2049_),
    .A2(_2051_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6214_ (.A1(_1405_),
    .A2(_3348_),
    .A3(_1947_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6215_ (.A1(_1946_),
    .A2(_2053_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6216_ (.I(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6217_ (.A1(_1882_),
    .A2(_1894_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6218_ (.A1(_1893_),
    .A2(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6219_ (.A1(_2057_),
    .A2(_1973_),
    .B(_1976_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6220_ (.A1(_1632_),
    .A2(_3378_),
    .A3(_1864_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6221_ (.A1(_1634_),
    .A2(_3362_),
    .A3(_1961_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6222_ (.A1(_1636_),
    .A2(_3362_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6223_ (.A1(_2059_),
    .A2(_2060_),
    .A3(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6224_ (.A1(_2059_),
    .A2(_2060_),
    .B(_2061_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6225_ (.A1(_2062_),
    .A2(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6226_ (.A1(_0358_),
    .A2(_3356_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6227_ (.A1(_2064_),
    .A2(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6228_ (.A1(_2058_),
    .A2(_2066_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6229_ (.A1(_2055_),
    .A2(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6230_ (.I(_1972_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6231_ (.A1(_1967_),
    .A2(_2069_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6232_ (.A1(_1967_),
    .A2(_1972_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6233_ (.A1(_1962_),
    .A2(_2071_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6234_ (.A1(_1981_),
    .A2(_1982_),
    .A3(_1987_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6235_ (.A1(_1980_),
    .A2(_2073_),
    .B(_1989_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6236_ (.A1(_1435_),
    .A2(_1039_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6237_ (.A1(_1437_),
    .A2(_3374_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6238_ (.A1(_1109_),
    .A2(\dspArea_regA[12] ),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6239_ (.A1(_2076_),
    .A2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6240_ (.A1(_2075_),
    .A2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6241_ (.A1(_0325_),
    .A2(_3390_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6242_ (.A1(_1443_),
    .A2(_3395_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6243_ (.A1(_1445_),
    .A2(_3403_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6244_ (.A1(_2081_),
    .A2(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6245_ (.A1(_2080_),
    .A2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6246_ (.A1(_1968_),
    .A2(_3398_),
    .A3(_1869_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6247_ (.A1(_1970_),
    .A2(_3385_),
    .A3(_1966_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6248_ (.A1(_2085_),
    .A2(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6249_ (.A1(_2079_),
    .A2(_2084_),
    .A3(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6250_ (.A1(_2074_),
    .A2(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6251_ (.A1(_2070_),
    .A2(_2072_),
    .A3(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6252_ (.A1(_2070_),
    .A2(_2072_),
    .B(_2089_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6253_ (.A1(_2090_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6254_ (.A1(_0829_),
    .A2(_3426_),
    .A3(_1889_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6255_ (.A1(_0608_),
    .A2(_3409_),
    .A3(_1986_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6256_ (.A1(_2093_),
    .A2(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6257_ (.A1(_0285_),
    .A2(_3450_),
    .A3(_1898_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6258_ (.A1(_0460_),
    .A2(_3434_),
    .A3(_1996_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6259_ (.A1(_0607_),
    .A2(_1884_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6260_ (.A1(_1234_),
    .A2(_3423_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6261_ (.A1(_1775_),
    .A2(_1992_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6262_ (.A1(_2099_),
    .A2(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6263_ (.A1(_2098_),
    .A2(_2101_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6264_ (.A1(_2096_),
    .A2(_2097_),
    .A3(_2102_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6265_ (.A1(_2096_),
    .A2(_2097_),
    .B(_2102_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6266_ (.A1(_2103_),
    .A2(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6267_ (.A1(_2095_),
    .A2(_2105_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6268_ (.A1(_0624_),
    .A2(_3440_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6269_ (.I(_3447_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6270_ (.A1(_0515_),
    .A2(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6271_ (.I(\dspArea_regA[21] ),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6272_ (.A1(_0468_),
    .A2(_2110_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6273_ (.A1(_2109_),
    .A2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6274_ (.A1(_2107_),
    .A2(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6275_ (.I(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6276_ (.A1(_1149_),
    .A2(_3465_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6277_ (.A1(_1367_),
    .A2(\dspArea_regA[23] ),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6278_ (.A1(\dspArea_regP[23] ),
    .A2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6279_ (.A1(_2115_),
    .A2(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6280_ (.A1(\dspArea_regP[22] ),
    .A2(_2000_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6281_ (.A1(_1999_),
    .A2(_2001_),
    .B(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6282_ (.A1(_2118_),
    .A2(_2120_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6283_ (.A1(_2114_),
    .A2(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6284_ (.A1(_2002_),
    .A2(_2004_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6285_ (.A1(_2002_),
    .A2(_2004_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6286_ (.A1(_1998_),
    .A2(_2123_),
    .B(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6287_ (.A1(_2122_),
    .A2(_2125_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6288_ (.A1(_2106_),
    .A2(_2126_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6289_ (.A1(_2005_),
    .A2(_2009_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6290_ (.A1(_1991_),
    .A2(_2010_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6291_ (.A1(_2128_),
    .A2(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6292_ (.A1(_2092_),
    .A2(_2127_),
    .A3(_2130_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6293_ (.A1(_2013_),
    .A2(_2014_),
    .A3(_2011_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6294_ (.A1(_2013_),
    .A2(_2014_),
    .B(_2011_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6295_ (.A1(_1977_),
    .A2(_2132_),
    .B(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6296_ (.A1(_2068_),
    .A2(_2131_),
    .A3(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6297_ (.A1(_2016_),
    .A2(_2019_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6298_ (.A1(_1951_),
    .A2(_2020_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6299_ (.A1(_2136_),
    .A2(_2137_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6300_ (.A1(_2052_),
    .A2(_2135_),
    .A3(_2138_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6301_ (.A1(_2048_),
    .A2(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6302_ (.A1(_2027_),
    .A2(_2030_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6303_ (.A1(_2027_),
    .A2(_2030_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6304_ (.A1(_2038_),
    .A2(_2040_),
    .B(_2142_),
    .C(_2141_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6305_ (.A1(_2141_),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6306_ (.A1(_2140_),
    .A2(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6307_ (.A1(_2140_),
    .A2(_2144_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6308_ (.A1(_2045_),
    .A2(_2145_),
    .A3(_2146_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6309_ (.A1(_3498_),
    .A2(_2044_),
    .A3(_2147_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6310_ (.A1(_2058_),
    .A2(_2066_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6311_ (.A1(_2055_),
    .A2(_2067_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6312_ (.A1(_2148_),
    .A2(_2149_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6313_ (.A1(_1405_),
    .A2(_3356_),
    .A3(_2064_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6314_ (.A1(_2063_),
    .A2(_2151_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6315_ (.I(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6316_ (.A1(_1980_),
    .A2(_1990_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6317_ (.A1(_1989_),
    .A2(_2154_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6318_ (.A1(_2155_),
    .A2(_2088_),
    .B(_2091_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6319_ (.A1(_1413_),
    .A2(_3386_),
    .A3(_1960_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6320_ (.A1(_1527_),
    .A2(_3370_),
    .A3(_2078_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6321_ (.A1(_1636_),
    .A2(_3370_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6322_ (.A1(_2157_),
    .A2(_2158_),
    .A3(_2159_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6323_ (.A1(_2157_),
    .A2(_2158_),
    .B(_2159_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6324_ (.A1(_2160_),
    .A2(_2161_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6325_ (.A1(_1533_),
    .A2(_3363_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6326_ (.A1(_2162_),
    .A2(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6327_ (.A1(_2156_),
    .A2(_2164_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6328_ (.A1(_2153_),
    .A2(_2165_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6329_ (.I(_2087_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6330_ (.A1(_2084_),
    .A2(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6331_ (.A1(_2084_),
    .A2(_2087_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6332_ (.A1(_2079_),
    .A2(_2169_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6333_ (.A1(_2096_),
    .A2(_2097_),
    .A3(_2102_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6334_ (.A1(_2095_),
    .A2(_2171_),
    .B(_2104_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6335_ (.A1(_1012_),
    .A2(_3376_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6336_ (.A1(_0995_),
    .A2(_3383_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6337_ (.A1(_0331_),
    .A2(_1058_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6338_ (.A1(_2174_),
    .A2(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6339_ (.A1(_2173_),
    .A2(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6340_ (.A1(_0747_),
    .A2(_3397_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6341_ (.A1(_0815_),
    .A2(_3404_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6342_ (.A1(_0313_),
    .A2(_3413_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6343_ (.A1(_2179_),
    .A2(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6344_ (.A1(_2178_),
    .A2(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6345_ (.A1(_1759_),
    .A2(_3407_),
    .A3(_1965_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6346_ (.A1(_0327_),
    .A2(_1346_),
    .A3(_2083_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6347_ (.A1(_2183_),
    .A2(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6348_ (.A1(_2177_),
    .A2(_2182_),
    .A3(_2185_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6349_ (.A1(_2172_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6350_ (.A1(_2168_),
    .A2(_2170_),
    .A3(_2187_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6351_ (.A1(_2168_),
    .A2(_2170_),
    .B(_2187_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6352_ (.A1(_2188_),
    .A2(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6353_ (.A1(_1225_),
    .A2(_3433_),
    .A3(_1985_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6354_ (.A1(_1342_),
    .A2(_1884_),
    .A3(_2101_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6355_ (.A1(_2191_),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6356_ (.A1(_1345_),
    .A2(_3458_),
    .A3(_1995_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6357_ (.A1(_1348_),
    .A2(_3442_),
    .A3(_2112_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6358_ (.A1(_1886_),
    .A2(_3424_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6359_ (.A1(_0604_),
    .A2(_1992_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6360_ (.A1(_1352_),
    .A2(_3438_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6361_ (.A1(_2197_),
    .A2(_2198_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6362_ (.A1(_2196_),
    .A2(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6363_ (.A1(_2194_),
    .A2(_2195_),
    .A3(_2200_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6364_ (.A1(_2194_),
    .A2(_2195_),
    .B(_2200_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6365_ (.A1(_2201_),
    .A2(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6366_ (.A1(_2193_),
    .A2(_2203_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6367_ (.A1(_0561_),
    .A2(_3448_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6368_ (.A1(_0282_),
    .A2(_2110_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6369_ (.A1(_0468_),
    .A2(\dspArea_regA[22] ),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6370_ (.A1(_2206_),
    .A2(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6371_ (.A1(_2205_),
    .A2(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6372_ (.I(_3472_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6373_ (.A1(_1150_),
    .A2(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6374_ (.A1(_0476_),
    .A2(\dspArea_regA[24] ),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6375_ (.A1(\dspArea_regP[24] ),
    .A2(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6376_ (.A1(_2211_),
    .A2(_2213_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6377_ (.A1(\dspArea_regP[23] ),
    .A2(_2116_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6378_ (.A1(_2115_),
    .A2(_2117_),
    .B(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6379_ (.A1(_2209_),
    .A2(_2214_),
    .A3(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6380_ (.A1(_2118_),
    .A2(_2120_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6381_ (.A1(_2118_),
    .A2(_2120_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6382_ (.A1(_2114_),
    .A2(_2218_),
    .B(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6383_ (.A1(_2217_),
    .A2(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6384_ (.A1(_2204_),
    .A2(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6385_ (.A1(_2122_),
    .A2(_2125_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6386_ (.A1(_2106_),
    .A2(_2126_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6387_ (.A1(_2223_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6388_ (.A1(_2190_),
    .A2(_2222_),
    .A3(_2225_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6389_ (.A1(_2128_),
    .A2(_2129_),
    .A3(_2127_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6390_ (.A1(_2128_),
    .A2(_2129_),
    .B(_2127_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6391_ (.A1(_2092_),
    .A2(_2227_),
    .B(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6392_ (.A1(_2166_),
    .A2(_2226_),
    .A3(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6393_ (.A1(_2131_),
    .A2(_2134_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6394_ (.A1(_2131_),
    .A2(_2134_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6395_ (.A1(_2068_),
    .A2(_2231_),
    .B(_2232_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6396_ (.A1(_2230_),
    .A2(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6397_ (.A1(_2150_),
    .A2(_2234_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6398_ (.A1(_2136_),
    .A2(_2137_),
    .A3(_2135_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6399_ (.A1(_2136_),
    .A2(_2137_),
    .B(_2135_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6400_ (.A1(_2052_),
    .A2(_2236_),
    .B(_2237_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6401_ (.A1(_2235_),
    .A2(_2238_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6402_ (.I(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6403_ (.A1(_2031_),
    .A2(_2140_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6404_ (.A1(_1821_),
    .A2(_1822_),
    .B(_2039_),
    .C(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6405_ (.A1(_2048_),
    .A2(_2139_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6406_ (.A1(_2141_),
    .A2(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6407_ (.A1(_2048_),
    .A2(_2139_),
    .B1(_2241_),
    .B2(_2037_),
    .C(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6408_ (.A1(_2242_),
    .A2(_2245_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6409_ (.A1(_1396_),
    .A2(_1504_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6410_ (.A1(_2247_),
    .A2(_1824_),
    .A3(_2039_),
    .A4(_2241_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6411_ (.A1(_1509_),
    .A2(_1510_),
    .B(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6412_ (.I(_2249_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6413_ (.A1(_2246_),
    .A2(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6414_ (.A1(_2240_),
    .A2(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6415_ (.I0(\dspArea_regP[24] ),
    .I1(_2252_),
    .S(_1619_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6416_ (.A1(_1932_),
    .A2(_2253_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6417_ (.I(\dspArea_regP[25] ),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6418_ (.A1(_2230_),
    .A2(_2233_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6419_ (.A1(_2150_),
    .A2(_2234_),
    .B(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6420_ (.A1(_2156_),
    .A2(_2164_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6421_ (.A1(_2153_),
    .A2(_2165_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6422_ (.A1(_2257_),
    .A2(_2258_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6423_ (.A1(_1407_),
    .A2(_3363_),
    .A3(_2162_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6424_ (.A1(_2161_),
    .A2(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6425_ (.A1(_2095_),
    .A2(_2105_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6426_ (.A1(_2104_),
    .A2(_2262_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6427_ (.A1(_2263_),
    .A2(_2186_),
    .B(_2189_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6428_ (.A1(_1414_),
    .A2(_3392_),
    .A3(_2077_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6429_ (.A1(_1845_),
    .A2(_3378_),
    .A3(_2176_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6430_ (.A1(_1847_),
    .A2(_3378_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6431_ (.A1(_2265_),
    .A2(_2266_),
    .A3(_2267_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6432_ (.A1(_2265_),
    .A2(_2266_),
    .B(_2267_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6433_ (.A1(_2268_),
    .A2(_2269_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6434_ (.A1(_0359_),
    .A2(_3371_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6435_ (.A1(_2270_),
    .A2(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6436_ (.A1(_2264_),
    .A2(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6437_ (.A1(_2261_),
    .A2(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6438_ (.I(_2185_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6439_ (.A1(_2182_),
    .A2(_2275_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6440_ (.A1(_2182_),
    .A2(_2185_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6441_ (.A1(_2177_),
    .A2(_2277_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6442_ (.A1(_2194_),
    .A2(_2195_),
    .A3(_2200_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6443_ (.A1(_2193_),
    .A2(_2279_),
    .B(_2202_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6444_ (.A1(_1435_),
    .A2(_3384_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6445_ (.A1(_1437_),
    .A2(_1058_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6446_ (.A1(_1323_),
    .A2(_1676_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6447_ (.A1(_2282_),
    .A2(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6448_ (.A1(_2281_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6449_ (.A1(_0927_),
    .A2(_3406_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6450_ (.A1(_1443_),
    .A2(_3413_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6451_ (.A1(_1445_),
    .A2(\dspArea_regA[17] ),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6452_ (.A1(_2287_),
    .A2(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6453_ (.A1(_2286_),
    .A2(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6454_ (.A1(_1968_),
    .A2(_3415_),
    .A3(_2082_),
    .Z(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6455_ (.A1(_1970_),
    .A2(_3398_),
    .A3(_2181_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6456_ (.A1(_2291_),
    .A2(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6457_ (.A1(_2285_),
    .A2(_2290_),
    .A3(_2293_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6458_ (.A1(_2280_),
    .A2(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6459_ (.A1(_2276_),
    .A2(_2278_),
    .A3(_2295_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6460_ (.A1(_2276_),
    .A2(_2278_),
    .B(_2295_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6461_ (.A1(_2296_),
    .A2(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6462_ (.A1(_0828_),
    .A2(_3441_),
    .A3(_2100_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6463_ (.A1(_0607_),
    .A2(_3425_),
    .A3(_2199_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6464_ (.A1(_2299_),
    .A2(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6465_ (.A1(_0547_),
    .A2(_3466_),
    .A3(_2111_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6466_ (.A1(_0562_),
    .A2(_3450_),
    .A3(_2208_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6467_ (.A1(_0306_),
    .A2(_3432_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6468_ (.A1(_1233_),
    .A2(_3438_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6469_ (.A1(_1134_),
    .A2(_3447_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6470_ (.A1(_2305_),
    .A2(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6471_ (.A1(_2304_),
    .A2(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6472_ (.A1(_2302_),
    .A2(_2303_),
    .A3(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6473_ (.A1(_2302_),
    .A2(_2303_),
    .B(_2308_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6474_ (.A1(_2309_),
    .A2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6475_ (.A1(_2301_),
    .A2(_2311_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6476_ (.A1(_0677_),
    .A2(_3457_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6477_ (.I(\dspArea_regA[22] ),
    .Z(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6478_ (.A1(_0464_),
    .A2(_2314_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6479_ (.A1(_0469_),
    .A2(\dspArea_regA[23] ),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6480_ (.A1(_2315_),
    .A2(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6481_ (.A1(_2313_),
    .A2(_2317_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6482_ (.I(\dspArea_regA[24] ),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6483_ (.A1(_1149_),
    .A2(_2319_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6484_ (.A1(_2254_),
    .A2(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6485_ (.A1(\dspArea_regP[24] ),
    .A2(_0265_),
    .A3(_2319_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6486_ (.I(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6487_ (.A1(_2211_),
    .A2(_2213_),
    .B(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6488_ (.A1(_2321_),
    .A2(_2324_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6489_ (.A1(_2318_),
    .A2(_2325_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6490_ (.I(_2209_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6491_ (.A1(_2214_),
    .A2(_2216_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6492_ (.A1(_2214_),
    .A2(_2216_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6493_ (.A1(_2327_),
    .A2(_2328_),
    .B(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6494_ (.A1(_2326_),
    .A2(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6495_ (.A1(_2312_),
    .A2(_2331_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6496_ (.A1(_2113_),
    .A2(_2121_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6497_ (.A1(_2219_),
    .A2(_2333_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6498_ (.A1(_2217_),
    .A2(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6499_ (.A1(_2204_),
    .A2(_2221_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6500_ (.A1(_2335_),
    .A2(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6501_ (.A1(_2298_),
    .A2(_2332_),
    .A3(_2337_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6502_ (.A1(_2223_),
    .A2(_2224_),
    .A3(_2222_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6503_ (.A1(_2223_),
    .A2(_2224_),
    .B(_2222_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6504_ (.A1(_2190_),
    .A2(_2339_),
    .B(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6505_ (.A1(_2338_),
    .A2(_2341_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6506_ (.A1(_2274_),
    .A2(_2342_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6507_ (.A1(_2226_),
    .A2(_2229_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6508_ (.A1(_2226_),
    .A2(_2229_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6509_ (.A1(_2166_),
    .A2(_2344_),
    .B(_2345_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6510_ (.A1(_2259_),
    .A2(_2343_),
    .A3(_2346_),
    .Z(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6511_ (.A1(_2256_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6512_ (.A1(_2235_),
    .A2(_2238_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6513_ (.A1(_2239_),
    .A2(_2251_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6514_ (.A1(_2349_),
    .A2(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6515_ (.A1(_2348_),
    .A2(_2351_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6516_ (.A1(_2045_),
    .A2(_2352_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6517_ (.I(_3490_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6518_ (.A1(_2254_),
    .A2(_0424_),
    .B(_2353_),
    .C(_2354_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6519_ (.I(\dspArea_regP[26] ),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6520_ (.A1(_2264_),
    .A2(_2272_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6521_ (.I(_2261_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6522_ (.A1(_2357_),
    .A2(_2273_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6523_ (.A1(_2356_),
    .A2(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6524_ (.A1(_1405_),
    .A2(_3371_),
    .A3(_2270_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6525_ (.A1(_2269_),
    .A2(_2360_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6526_ (.I(_2361_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6527_ (.A1(_2193_),
    .A2(_2203_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6528_ (.A1(_2202_),
    .A2(_2363_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6529_ (.A1(_2364_),
    .A2(_2294_),
    .B(_2297_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6530_ (.A1(_1632_),
    .A2(_3400_),
    .A3(_2175_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6531_ (.A1(_1527_),
    .A2(_3386_),
    .A3(_2284_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6532_ (.A1(_1636_),
    .A2(_3386_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6533_ (.A1(_2366_),
    .A2(_2367_),
    .A3(_2368_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6534_ (.A1(_2366_),
    .A2(_2367_),
    .B(_2368_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6535_ (.A1(_2369_),
    .A2(_2370_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6536_ (.A1(_1533_),
    .A2(_3379_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6537_ (.A1(_2371_),
    .A2(_2372_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6538_ (.A1(_2365_),
    .A2(_2373_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6539_ (.A1(_2362_),
    .A2(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6540_ (.I(_2293_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6541_ (.A1(_2290_),
    .A2(_2376_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6542_ (.A1(_2290_),
    .A2(_2293_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6543_ (.A1(_2285_),
    .A2(_2378_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6544_ (.A1(_2302_),
    .A2(_2303_),
    .A3(_2308_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6545_ (.A1(_2301_),
    .A2(_2380_),
    .B(_2310_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6546_ (.A1(_1011_),
    .A2(_1059_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6547_ (.A1(\dspArea_regB[12] ),
    .A2(_1676_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6548_ (.A1(_0330_),
    .A2(\dspArea_regA[15] ),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6549_ (.A1(_2383_),
    .A2(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6550_ (.A1(_2382_),
    .A2(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6551_ (.A1(_0926_),
    .A2(_3414_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6552_ (.A1(_0318_),
    .A2(\dspArea_regA[17] ),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6553_ (.A1(_0312_),
    .A2(\dspArea_regA[18] ),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6554_ (.A1(_2388_),
    .A2(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6555_ (.A1(_2387_),
    .A2(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6556_ (.A1(_0321_),
    .A2(_1582_),
    .A3(_2180_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6557_ (.A1(_0326_),
    .A2(_3406_),
    .A3(_2289_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6558_ (.A1(_2392_),
    .A2(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6559_ (.A1(_2386_),
    .A2(_2391_),
    .A3(_2394_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6560_ (.A1(_2381_),
    .A2(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6561_ (.A1(_2377_),
    .A2(_2379_),
    .A3(_2396_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6562_ (.A1(_2377_),
    .A2(_2379_),
    .B(_2396_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6563_ (.A1(_2397_),
    .A2(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6564_ (.A1(_0828_),
    .A2(_3450_),
    .A3(_2198_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6565_ (.A1(_0760_),
    .A2(_3433_),
    .A3(_2307_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6566_ (.A1(_2400_),
    .A2(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6567_ (.A1(_0464_),
    .A2(_3472_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6568_ (.I(_2403_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6569_ (.A1(_2207_),
    .A2(_2404_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6570_ (.A1(_0562_),
    .A2(_3458_),
    .A3(_2317_),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6571_ (.A1(_0614_),
    .A2(_3440_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6572_ (.A1(_1233_),
    .A2(_2108_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6573_ (.A1(_1134_),
    .A2(\dspArea_regA[21] ),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6574_ (.A1(_2408_),
    .A2(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6575_ (.A1(_2407_),
    .A2(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6576_ (.A1(_2405_),
    .A2(_2406_),
    .A3(_2411_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6577_ (.A1(_2405_),
    .A2(_2406_),
    .B(_2411_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6578_ (.A1(_2412_),
    .A2(_2413_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6579_ (.A1(_2402_),
    .A2(_2414_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6580_ (.A1(\dspArea_regP[25] ),
    .A2(_1150_),
    .A3(_3478_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6581_ (.A1(\dspArea_regP[26] ),
    .A2(_2416_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6582_ (.A1(_0622_),
    .A2(_2314_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6583_ (.A1(_0278_),
    .A2(_3478_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6584_ (.A1(_2403_),
    .A2(_2418_),
    .A3(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6585_ (.A1(_2417_),
    .A2(_2420_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6586_ (.A1(_2321_),
    .A2(_2324_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6587_ (.A1(_2318_),
    .A2(_2325_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6588_ (.A1(_2422_),
    .A2(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6589_ (.A1(_2415_),
    .A2(_2421_),
    .A3(_2424_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6590_ (.A1(_2326_),
    .A2(_2330_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6591_ (.A1(_2312_),
    .A2(_2331_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6592_ (.A1(_2426_),
    .A2(_2427_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6593_ (.A1(_2399_),
    .A2(_2425_),
    .A3(_2428_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6594_ (.A1(_2335_),
    .A2(_2336_),
    .A3(_2332_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6595_ (.A1(_2335_),
    .A2(_2336_),
    .B(_2332_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6596_ (.A1(_2298_),
    .A2(_2430_),
    .B(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6597_ (.A1(_2375_),
    .A2(_2429_),
    .A3(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6598_ (.A1(_2338_),
    .A2(_2341_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6599_ (.A1(_2274_),
    .A2(_2342_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6600_ (.A1(_2434_),
    .A2(_2435_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6601_ (.A1(_2359_),
    .A2(_2433_),
    .A3(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6602_ (.A1(_2343_),
    .A2(_2346_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6603_ (.A1(_2343_),
    .A2(_2346_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6604_ (.A1(_2259_),
    .A2(_2438_),
    .B(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6605_ (.A1(_2437_),
    .A2(_2440_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6606_ (.A1(_2259_),
    .A2(_2438_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6607_ (.A1(_2259_),
    .A2(_2438_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6608_ (.A1(_2256_),
    .A2(_2442_),
    .A3(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6609_ (.A1(_2150_),
    .A2(_2234_),
    .B(_2347_),
    .C(_2255_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6610_ (.A1(_2235_),
    .A2(_2238_),
    .A3(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6611_ (.A1(_2444_),
    .A2(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6612_ (.I(_2348_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6613_ (.A1(_2246_),
    .A2(_2250_),
    .B(_2448_),
    .C(_2240_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6614_ (.A1(_2441_),
    .A2(_2447_),
    .A3(_2449_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6615_ (.A1(_2447_),
    .A2(_2449_),
    .B(_2441_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6616_ (.A1(_2450_),
    .A2(_2451_),
    .B(_0367_),
    .C(_0986_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6617_ (.A1(_2355_),
    .A2(_0424_),
    .B(_2452_),
    .C(_2354_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6618_ (.I(\dspArea_regP[27] ),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6619_ (.I(_0422_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6620_ (.A1(_2434_),
    .A2(_2435_),
    .A3(_2433_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6621_ (.A1(_2434_),
    .A2(_2435_),
    .B(_2433_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6622_ (.A1(_2359_),
    .A2(_2455_),
    .B(_2456_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6623_ (.A1(_2365_),
    .A2(_2373_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6624_ (.A1(_2362_),
    .A2(_2374_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6625_ (.A1(_2458_),
    .A2(_2459_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6626_ (.A1(_1297_),
    .A2(_3379_),
    .A3(_2371_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6627_ (.A1(_2370_),
    .A2(_2461_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6628_ (.I(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6629_ (.A1(_2301_),
    .A2(_2311_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6630_ (.A1(_2310_),
    .A2(_2464_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6631_ (.A1(_2465_),
    .A2(_2395_),
    .B(_2398_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6632_ (.A1(\dspArea_regB[12] ),
    .A2(_3403_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6633_ (.A1(_2283_),
    .A2(_2467_),
    .Z(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6634_ (.A1(_1305_),
    .A2(_3392_),
    .A3(_2385_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6635_ (.A1(_0352_),
    .A2(_3392_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6636_ (.A1(_2468_),
    .A2(_2469_),
    .A3(_2470_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6637_ (.A1(_2468_),
    .A2(_2469_),
    .B(_2470_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6638_ (.A1(_2471_),
    .A2(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6639_ (.A1(_1197_),
    .A2(_3387_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6640_ (.A1(_2473_),
    .A2(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6641_ (.A1(_2466_),
    .A2(_2475_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6642_ (.A1(_2463_),
    .A2(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6643_ (.I(_2394_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6644_ (.A1(_2391_),
    .A2(_2478_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6645_ (.A1(_2391_),
    .A2(_2394_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6646_ (.A1(_2386_),
    .A2(_2480_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6647_ (.A1(_2405_),
    .A2(_2406_),
    .A3(_2411_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6648_ (.A1(_2402_),
    .A2(_2482_),
    .B(_2413_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6649_ (.A1(_1011_),
    .A2(_3396_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6650_ (.A1(_1323_),
    .A2(_1368_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6651_ (.A1(_2467_),
    .A2(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6652_ (.A1(_2484_),
    .A2(_2486_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6653_ (.A1(_1018_),
    .A2(_3423_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6654_ (.A1(_0735_),
    .A2(\dspArea_regA[18] ),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6655_ (.A1(_1116_),
    .A2(\dspArea_regA[19] ),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6656_ (.A1(_2489_),
    .A2(_2490_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6657_ (.A1(_2488_),
    .A2(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6658_ (.I(_3432_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6659_ (.A1(_0924_),
    .A2(_2493_),
    .A3(_2288_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6660_ (.A1(_1450_),
    .A2(_3415_),
    .A3(_2390_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6661_ (.A1(_2494_),
    .A2(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6662_ (.A1(_2487_),
    .A2(_2492_),
    .A3(_2496_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6663_ (.A1(_2483_),
    .A2(_2497_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6664_ (.A1(_2479_),
    .A2(_2481_),
    .A3(_2498_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6665_ (.A1(_2479_),
    .A2(_2481_),
    .B(_2498_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6666_ (.A1(_2499_),
    .A2(_2500_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6667_ (.A1(_0284_),
    .A2(_3479_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6668_ (.A1(_0624_),
    .A2(_2210_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6669_ (.A1(_2502_),
    .A2(_2503_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6670_ (.A1(_0561_),
    .A2(_3478_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6671_ (.A1(_2404_),
    .A2(_2505_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6672_ (.A1(_2504_),
    .A2(_2506_),
    .B(_2453_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6673_ (.A1(_2453_),
    .A2(_2504_),
    .A3(_2506_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6674_ (.A1(_2507_),
    .A2(_2508_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6675_ (.A1(\dspArea_regP[26] ),
    .A2(_2416_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6676_ (.A1(_2417_),
    .A2(_2420_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6677_ (.A1(_2510_),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6678_ (.A1(_2509_),
    .A2(_2512_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6679_ (.A1(_1233_),
    .A2(_2110_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6680_ (.A1(_2306_),
    .A2(_2514_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6681_ (.A1(_0760_),
    .A2(_3442_),
    .A3(_2410_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6682_ (.A1(_2515_),
    .A2(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6683_ (.I(_2418_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6684_ (.A1(_2404_),
    .A2(_2419_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6685_ (.A1(_0279_),
    .A2(_3479_),
    .A3(_2404_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6686_ (.A1(_2518_),
    .A2(_2519_),
    .B(_2520_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6687_ (.A1(\dspArea_regB[7] ),
    .A2(_2108_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6688_ (.A1(_1775_),
    .A2(_3465_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6689_ (.A1(_2514_),
    .A2(_2522_),
    .A3(_2523_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6690_ (.A1(_2521_),
    .A2(_2524_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6691_ (.A1(_2517_),
    .A2(_2525_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6692_ (.A1(_2513_),
    .A2(_2526_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6693_ (.A1(_2422_),
    .A2(_2423_),
    .A3(_2421_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6694_ (.A1(_2422_),
    .A2(_2423_),
    .B(_2421_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6695_ (.A1(_2415_),
    .A2(_2528_),
    .B(_2529_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6696_ (.A1(_2527_),
    .A2(_2530_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6697_ (.A1(_2501_),
    .A2(_2531_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6698_ (.A1(_2426_),
    .A2(_2427_),
    .A3(_2425_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6699_ (.A1(_2426_),
    .A2(_2427_),
    .B(_2425_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6700_ (.A1(_2399_),
    .A2(_2533_),
    .B(_2534_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6701_ (.A1(_2477_),
    .A2(_2532_),
    .A3(_2535_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6702_ (.A1(_2429_),
    .A2(_2432_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6703_ (.A1(_2429_),
    .A2(_2432_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6704_ (.A1(_2375_),
    .A2(_2537_),
    .B(_2538_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6705_ (.A1(_2536_),
    .A2(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6706_ (.A1(_2460_),
    .A2(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6707_ (.A1(_2457_),
    .A2(_2541_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6708_ (.A1(_2437_),
    .A2(_2440_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6709_ (.A1(_2543_),
    .A2(_2451_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6710_ (.A1(_2542_),
    .A2(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6711_ (.A1(_2542_),
    .A2(_2544_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6712_ (.A1(_0423_),
    .A2(_2545_),
    .A3(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6713_ (.A1(_2453_),
    .A2(_2454_),
    .B(_2547_),
    .C(_2354_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6714_ (.A1(_2466_),
    .A2(_2475_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6715_ (.A1(_2463_),
    .A2(_2476_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6716_ (.A1(_2548_),
    .A2(_2549_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6717_ (.A1(_1519_),
    .A2(_3387_),
    .A3(_2473_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6718_ (.A1(_2472_),
    .A2(_2551_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6719_ (.I(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6720_ (.A1(_2402_),
    .A2(_2414_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6721_ (.A1(_2413_),
    .A2(_2554_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6722_ (.A1(_2555_),
    .A2(_2497_),
    .B(_2500_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6723_ (.A1(_0334_),
    .A2(_3416_),
    .A3(_2467_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6724_ (.A1(_1527_),
    .A2(_3400_),
    .A3(_2486_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6725_ (.A1(_1418_),
    .A2(_3400_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6726_ (.A1(_2557_),
    .A2(_2558_),
    .A3(_2559_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6727_ (.A1(_2557_),
    .A2(_2558_),
    .B(_2559_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6728_ (.A1(_2560_),
    .A2(_2561_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6729_ (.A1(_1533_),
    .A2(_3393_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6730_ (.A1(_2562_),
    .A2(_2563_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6731_ (.A1(_2556_),
    .A2(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6732_ (.A1(_2553_),
    .A2(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6733_ (.A1(\dspArea_regP[28] ),
    .A2(_2505_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6734_ (.A1(_2514_),
    .A2(_2523_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6735_ (.A1(_0604_),
    .A2(_2314_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6736_ (.A1(_2409_),
    .A2(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6737_ (.A1(_2522_),
    .A2(_2568_),
    .B(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6738_ (.A1(_0305_),
    .A2(_3456_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6739_ (.A1(_0297_),
    .A2(_2210_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6740_ (.A1(_2569_),
    .A2(_2572_),
    .A3(_2573_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6741_ (.A1(_2506_),
    .A2(_2574_),
    .Z(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6742_ (.A1(_2571_),
    .A2(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6743_ (.A1(_2508_),
    .A2(_2567_),
    .A3(_2576_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6744_ (.A1(_2510_),
    .A2(_2511_),
    .B(_2509_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6745_ (.I(_2578_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6746_ (.A1(_2513_),
    .A2(_2526_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6747_ (.A1(_2579_),
    .A2(_2580_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6748_ (.A1(_2494_),
    .A2(_2495_),
    .B(_2492_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6749_ (.A1(_2494_),
    .A2(_2495_),
    .A3(_2492_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6750_ (.A1(_2487_),
    .A2(_2583_),
    .A3(_2582_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6751_ (.A1(_2582_),
    .A2(_2584_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6752_ (.A1(_2521_),
    .A2(_2524_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6753_ (.I(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6754_ (.A1(_2517_),
    .A2(_2525_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6755_ (.A1(_2587_),
    .A2(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6756_ (.A1(_1013_),
    .A2(_3407_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6757_ (.A1(_0341_),
    .A2(_1478_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6758_ (.A1(_0332_),
    .A2(_1582_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6759_ (.A1(_2591_),
    .A2(_2592_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6760_ (.A1(_2590_),
    .A2(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6761_ (.A1(_1968_),
    .A2(_3441_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6762_ (.A1(_1450_),
    .A2(_2493_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6763_ (.A1(_0314_),
    .A2(_3449_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6764_ (.A1(_2595_),
    .A2(_2596_),
    .A3(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6765_ (.A1(_0323_),
    .A2(_3443_),
    .A3(_2389_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6766_ (.A1(_0748_),
    .A2(_3426_),
    .A3(_2491_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6767_ (.A1(_2599_),
    .A2(_2600_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6768_ (.A1(_2594_),
    .A2(_2598_),
    .A3(_2601_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6769_ (.A1(_2585_),
    .A2(_2589_),
    .A3(_2602_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6770_ (.A1(_2577_),
    .A2(_2581_),
    .A3(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6771_ (.I(_2527_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6772_ (.A1(_2605_),
    .A2(_2530_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6773_ (.A1(_2501_),
    .A2(_2531_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6774_ (.A1(_2606_),
    .A2(_2607_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6775_ (.A1(_2566_),
    .A2(_2604_),
    .A3(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6776_ (.A1(_2532_),
    .A2(_2535_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6777_ (.A1(_2532_),
    .A2(_2535_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6778_ (.A1(_2477_),
    .A2(_2610_),
    .B(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6779_ (.A1(_2609_),
    .A2(_2612_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6780_ (.A1(_2536_),
    .A2(_2539_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6781_ (.A1(_2460_),
    .A2(_2540_),
    .B(_2614_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6782_ (.A1(_2550_),
    .A2(_2613_),
    .A3(_2615_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6783_ (.A1(_2457_),
    .A2(_2541_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6784_ (.A1(_2437_),
    .A2(_2440_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6785_ (.A1(_2444_),
    .A2(_2446_),
    .B(_2617_),
    .C(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6786_ (.A1(_2457_),
    .A2(_2541_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6787_ (.A1(_2457_),
    .A2(_2541_),
    .B(_2437_),
    .C(_2440_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6788_ (.A1(_2620_),
    .A2(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6789_ (.A1(_2239_),
    .A2(_2348_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6790_ (.A1(_2441_),
    .A2(_2542_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6791_ (.A1(_2246_),
    .A2(_2250_),
    .B(_2623_),
    .C(_2624_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6792_ (.A1(_2619_),
    .A2(_2622_),
    .A3(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6793_ (.A1(_2616_),
    .A2(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6794_ (.I(_0395_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6795_ (.I0(\dspArea_regP[28] ),
    .I1(_2627_),
    .S(_2628_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6796_ (.A1(_1932_),
    .A2(_2629_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6797_ (.I(_2550_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6798_ (.I(_2613_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6799_ (.A1(_2609_),
    .A2(_2612_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6800_ (.A1(_2630_),
    .A2(_2631_),
    .B(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6801_ (.A1(_2556_),
    .A2(_2564_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6802_ (.A1(_2553_),
    .A2(_2565_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6803_ (.A1(_2634_),
    .A2(_2635_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6804_ (.A1(\dspArea_regP[28] ),
    .A2(_2505_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6805_ (.A1(\dspArea_regP[29] ),
    .A2(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6806_ (.A1(_1886_),
    .A2(_3466_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6807_ (.A1(_0839_),
    .A2(_3472_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6808_ (.A1(_1775_),
    .A2(_2319_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6809_ (.A1(_2640_),
    .A2(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6810_ (.A1(_2639_),
    .A2(_2642_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6811_ (.A1(_2569_),
    .A2(_2573_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6812_ (.A1(_2523_),
    .A2(_2640_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6813_ (.A1(_2572_),
    .A2(_2644_),
    .B(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6814_ (.A1(_2643_),
    .A2(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6815_ (.A1(_2638_),
    .A2(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6816_ (.A1(_2508_),
    .A2(_2567_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6817_ (.A1(_2508_),
    .A2(_2567_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6818_ (.A1(_2649_),
    .A2(_2576_),
    .B(_2650_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6819_ (.A1(_2648_),
    .A2(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6820_ (.A1(_2599_),
    .A2(_2600_),
    .A3(_2598_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6821_ (.A1(_2599_),
    .A2(_2600_),
    .B(_2598_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6822_ (.A1(_2594_),
    .A2(_2653_),
    .B(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6823_ (.A1(_2506_),
    .A2(_2574_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6824_ (.A1(_2571_),
    .A2(_2575_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6825_ (.A1(_2656_),
    .A2(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6826_ (.A1(_1305_),
    .A2(_3416_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6827_ (.A1(_0341_),
    .A2(_3424_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6828_ (.A1(_0333_),
    .A2(_2493_),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6829_ (.A1(_2660_),
    .A2(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6830_ (.A1(_2659_),
    .A2(_2662_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6831_ (.A1(_0928_),
    .A2(_3440_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6832_ (.A1(_0736_),
    .A2(_3448_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6833_ (.A1(_1755_),
    .A2(_3456_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6834_ (.A1(_2665_),
    .A2(_2666_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6835_ (.A1(_2664_),
    .A2(_2667_),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6836_ (.A1(_2595_),
    .A2(_2597_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6837_ (.A1(_2490_),
    .A2(_2665_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6838_ (.A1(_2596_),
    .A2(_2669_),
    .B(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6839_ (.A1(_2668_),
    .A2(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6840_ (.A1(_2663_),
    .A2(_2672_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6841_ (.A1(_2655_),
    .A2(_2658_),
    .A3(_2673_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6842_ (.A1(_2652_),
    .A2(_2674_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6843_ (.I(_2675_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6844_ (.A1(_2579_),
    .A2(_2580_),
    .A3(_2577_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6845_ (.A1(_2579_),
    .A2(_2580_),
    .B(_2577_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6846_ (.A1(_2677_),
    .A2(_2603_),
    .B(_2678_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6847_ (.A1(_0361_),
    .A2(_3393_),
    .A3(_2562_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6848_ (.A1(_2561_),
    .A2(_2680_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6849_ (.A1(_2587_),
    .A2(_2588_),
    .A3(_2602_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6850_ (.A1(_2587_),
    .A2(_2588_),
    .B(_2602_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6851_ (.A1(_2585_),
    .A2(_2682_),
    .B(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6852_ (.A1(_2590_),
    .A2(_2593_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6853_ (.A1(_2485_),
    .A2(_2660_),
    .B(_2685_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6854_ (.A1(_0353_),
    .A2(_3409_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6855_ (.A1(_2686_),
    .A2(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6856_ (.A1(_1198_),
    .A2(_3401_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6857_ (.A1(_2688_),
    .A2(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6858_ (.A1(_2684_),
    .A2(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6859_ (.A1(_2681_),
    .A2(_2691_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6860_ (.A1(_2676_),
    .A2(_2679_),
    .A3(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6861_ (.A1(_2606_),
    .A2(_2607_),
    .A3(_2604_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6862_ (.A1(_2606_),
    .A2(_2607_),
    .B(_2604_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6863_ (.A1(_2566_),
    .A2(_2694_),
    .B(_2695_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6864_ (.A1(_2636_),
    .A2(_2693_),
    .A3(_2696_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6865_ (.A1(_2633_),
    .A2(_2697_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6866_ (.I(_2616_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6867_ (.A1(_2630_),
    .A2(_2631_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6868_ (.A1(_2630_),
    .A2(_2631_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6869_ (.A1(_2700_),
    .A2(_2701_),
    .A3(_2615_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6870_ (.A1(_2699_),
    .A2(_2626_),
    .B(_2702_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6871_ (.A1(_2698_),
    .A2(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6872_ (.A1(\dspArea_regP[29] ),
    .A2(_0380_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6873_ (.A1(_0988_),
    .A2(_2704_),
    .B(_2705_),
    .C(_2354_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6874_ (.A1(_0828_),
    .A2(_3480_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6875_ (.A1(_0760_),
    .A2(_3473_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6876_ (.A1(_2706_),
    .A2(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6877_ (.A1(_2706_),
    .A2(_2707_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6878_ (.A1(_2708_),
    .A2(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6879_ (.A1(_0298_),
    .A2(_3480_),
    .A3(_2640_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6880_ (.A1(_2639_),
    .A2(_2642_),
    .B(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6881_ (.A1(_2710_),
    .A2(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6882_ (.A1(\dspArea_regP[30] ),
    .A2(_2713_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6883_ (.A1(\dspArea_regP[29] ),
    .A2(_2637_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6884_ (.A1(_2638_),
    .A2(_2647_),
    .B(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6885_ (.A1(_2714_),
    .A2(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6886_ (.I(_2663_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6887_ (.A1(_2668_),
    .A2(_2671_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6888_ (.A1(_2718_),
    .A2(_2672_),
    .B(_2719_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6889_ (.A1(_2643_),
    .A2(_2646_),
    .Z(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6890_ (.A1(_0347_),
    .A2(_3424_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6891_ (.A1(_0996_),
    .A2(_1992_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6892_ (.A1(_1110_),
    .A2(_3439_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6893_ (.A1(_2723_),
    .A2(_2724_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6894_ (.A1(_2722_),
    .A2(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6895_ (.A1(_0928_),
    .A2(_3449_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6896_ (.A1(_0736_),
    .A2(_2110_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6897_ (.A1(_1755_),
    .A2(_2314_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6898_ (.A1(_2728_),
    .A2(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6899_ (.A1(_2727_),
    .A2(_2730_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6900_ (.A1(_0323_),
    .A2(_3459_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6901_ (.A1(_2597_),
    .A2(_2732_),
    .B1(_2667_),
    .B2(_2664_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6902_ (.A1(_2726_),
    .A2(_2731_),
    .A3(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6903_ (.A1(_2721_),
    .A2(_2734_),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6904_ (.A1(_2720_),
    .A2(_2735_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6905_ (.A1(_2717_),
    .A2(_2736_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6906_ (.A1(_2638_),
    .A2(_2647_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6907_ (.A1(_2638_),
    .A2(_2647_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6908_ (.A1(_2738_),
    .A2(_2739_),
    .A3(_2651_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6909_ (.A1(_2652_),
    .A2(_2674_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6910_ (.A1(_2740_),
    .A2(_2741_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6911_ (.A1(_2737_),
    .A2(_2742_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6912_ (.A1(_0356_),
    .A2(_3410_),
    .A3(_2686_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6913_ (.A1(_0361_),
    .A2(_3401_),
    .A3(_2688_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6914_ (.A1(_2744_),
    .A2(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6915_ (.I(_2655_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6916_ (.A1(_2658_),
    .A2(_2673_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6917_ (.A1(_2658_),
    .A2(_2673_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6918_ (.A1(_2747_),
    .A2(_2748_),
    .B(_2749_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6919_ (.A1(_1632_),
    .A2(_3434_),
    .A3(_2592_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6920_ (.A1(_0349_),
    .A2(_3416_),
    .A3(_2662_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6921_ (.A1(_2751_),
    .A2(_2752_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6922_ (.A1(_1419_),
    .A2(_3417_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6923_ (.A1(_2753_),
    .A2(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6924_ (.A1(_1424_),
    .A2(_3409_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6925_ (.A1(_2755_),
    .A2(_2756_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6926_ (.A1(_2750_),
    .A2(_2757_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6927_ (.A1(_2746_),
    .A2(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6928_ (.A1(_2676_),
    .A2(_2679_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6929_ (.A1(_2676_),
    .A2(_2679_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6930_ (.A1(_2760_),
    .A2(_2692_),
    .B(_2761_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6931_ (.A1(_2743_),
    .A2(_2759_),
    .A3(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6932_ (.A1(_2684_),
    .A2(_2690_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6933_ (.A1(_2681_),
    .A2(_2691_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6934_ (.A1(_2764_),
    .A2(_2765_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6935_ (.A1(_2763_),
    .A2(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6936_ (.A1(_2693_),
    .A2(_2696_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6937_ (.A1(_2693_),
    .A2(_2696_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6938_ (.A1(_2636_),
    .A2(_2768_),
    .B(_2769_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6939_ (.A1(_2767_),
    .A2(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6940_ (.A1(_2636_),
    .A2(_2768_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6941_ (.A1(_2636_),
    .A2(_2768_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6942_ (.A1(_2633_),
    .A2(_2772_),
    .A3(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6943_ (.A1(_2630_),
    .A2(_2631_),
    .B(_2697_),
    .C(_2632_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6944_ (.A1(_2700_),
    .A2(_2701_),
    .A3(_2615_),
    .A4(_2775_),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6945_ (.A1(_2774_),
    .A2(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6946_ (.A1(_2616_),
    .A2(_2698_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6947_ (.I(_2778_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6948_ (.A1(_2619_),
    .A2(_2622_),
    .A3(_2625_),
    .B(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6949_ (.A1(_2777_),
    .A2(_2780_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6950_ (.A1(_2771_),
    .A2(_2781_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6951_ (.I0(\dspArea_regP[30] ),
    .I1(_2782_),
    .S(_2628_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6952_ (.A1(_1932_),
    .A2(_2783_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6953_ (.I(\dspArea_regP[31] ),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6954_ (.I(_2767_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6955_ (.A1(_2785_),
    .A2(_2770_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6956_ (.A1(_2785_),
    .A2(_2770_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6957_ (.A1(_2777_),
    .A2(_2780_),
    .B(_2787_),
    .C(_2786_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6958_ (.A1(_2743_),
    .A2(_2759_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6959_ (.A1(_2743_),
    .A2(_2759_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6960_ (.A1(_2789_),
    .A2(_2790_),
    .A3(_2762_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6961_ (.A1(_2763_),
    .A2(_2766_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6962_ (.A1(\dspArea_regP[30] ),
    .A2(_2713_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6963_ (.I(_0309_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6964_ (.I(_3481_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6965_ (.A1(_2794_),
    .A2(_2795_),
    .A3(_2640_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6966_ (.A1(\dspArea_regP[31] ),
    .A2(_2796_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6967_ (.A1(_2793_),
    .A2(_2797_),
    .Z(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6968_ (.I(_2726_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6969_ (.A1(_2731_),
    .A2(_2733_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6970_ (.A1(_2731_),
    .A2(_2733_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6971_ (.A1(_2799_),
    .A2(_2800_),
    .B(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6972_ (.A1(_2708_),
    .A2(_2709_),
    .A3(_2712_),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6973_ (.A1(_0347_),
    .A2(_2493_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6974_ (.A1(_0996_),
    .A2(_3439_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6975_ (.A1(_1110_),
    .A2(_2108_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6976_ (.A1(_2805_),
    .A2(_2806_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6977_ (.A1(_2804_),
    .A2(_2807_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6978_ (.A1(_1970_),
    .A2(_3457_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6979_ (.A1(_0320_),
    .A2(_3465_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6980_ (.A1(_1755_),
    .A2(\dspArea_regA[23] ),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6981_ (.A1(_2810_),
    .A2(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6982_ (.A1(_2809_),
    .A2(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6983_ (.A1(_0315_),
    .A2(_3467_),
    .A3(_2728_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6984_ (.A1(_2727_),
    .A2(_2730_),
    .B(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6985_ (.A1(_2808_),
    .A2(_2813_),
    .A3(_2815_),
    .Z(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6986_ (.A1(_2803_),
    .A2(_2816_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6987_ (.A1(_2802_),
    .A2(_2817_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6988_ (.A1(_2798_),
    .A2(_2818_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6989_ (.A1(_2714_),
    .A2(_2716_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6990_ (.A1(_2717_),
    .A2(_2736_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6991_ (.A1(_2820_),
    .A2(_2821_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6992_ (.A1(_2819_),
    .A2(_2822_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6993_ (.I(_2753_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6994_ (.A1(_2824_),
    .A2(_2754_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6995_ (.A1(_0361_),
    .A2(_3410_),
    .A3(_2755_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6996_ (.A1(_2825_),
    .A2(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6997_ (.A1(_2721_),
    .A2(_2734_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6998_ (.A1(_2720_),
    .A2(_2735_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6999_ (.A1(_2828_),
    .A2(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7000_ (.A1(_1190_),
    .A2(_3443_),
    .A3(_2661_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7001_ (.A1(_0349_),
    .A2(_3426_),
    .A3(_2725_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7002_ (.A1(_2831_),
    .A2(_2832_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7003_ (.A1(_1419_),
    .A2(_3427_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7004_ (.A1(_2833_),
    .A2(_2834_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7005_ (.A1(_1424_),
    .A2(_3417_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7006_ (.A1(_2835_),
    .A2(_2836_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7007_ (.A1(_2830_),
    .A2(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7008_ (.A1(_2827_),
    .A2(_2838_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7009_ (.A1(_2823_),
    .A2(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7010_ (.I(_2737_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7011_ (.A1(_2841_),
    .A2(_2742_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7012_ (.A1(_2842_),
    .A2(_2790_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7013_ (.A1(_2750_),
    .A2(_2757_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7014_ (.A1(_2744_),
    .A2(_2745_),
    .B(_2758_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7015_ (.A1(_2844_),
    .A2(_2845_),
    .Z(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _7016_ (.A1(_2840_),
    .A2(_2843_),
    .A3(_2846_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7017_ (.A1(_2791_),
    .A2(_2792_),
    .A3(_2847_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7018_ (.A1(_2791_),
    .A2(_2792_),
    .B(_2847_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7019_ (.A1(_2848_),
    .A2(_2849_),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7020_ (.I(_2850_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7021_ (.A1(_2786_),
    .A2(_2788_),
    .A3(_2851_),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7022_ (.A1(_2786_),
    .A2(_2788_),
    .B(_2851_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7023_ (.A1(_1831_),
    .A2(_2852_),
    .A3(_2853_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7024_ (.I(_3490_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7025_ (.A1(_2784_),
    .A2(_2454_),
    .B(_2854_),
    .C(_2855_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7026_ (.I(_3558_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7027_ (.A1(\dspArea_regP[31] ),
    .A2(_2796_),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7028_ (.A1(\dspArea_regP[32] ),
    .A2(_2857_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7029_ (.A1(_2706_),
    .A2(_2707_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7030_ (.I(_2808_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7031_ (.A1(_2813_),
    .A2(_2815_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7032_ (.A1(_2813_),
    .A2(_2815_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7033_ (.A1(_2860_),
    .A2(_2861_),
    .B(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7034_ (.A1(_0348_),
    .A2(_3441_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7035_ (.A1(_0996_),
    .A2(_3449_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7036_ (.A1(_0332_),
    .A2(_3457_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7037_ (.A1(_2865_),
    .A2(_2866_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7038_ (.A1(_2864_),
    .A2(_2867_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7039_ (.A1(_0737_),
    .A2(_2210_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7040_ (.A1(_0314_),
    .A2(_2319_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7041_ (.A1(_2869_),
    .A2(_2870_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7042_ (.A1(_0327_),
    .A2(_3467_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7043_ (.A1(_2871_),
    .A2(_2872_),
    .Z(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7044_ (.A1(_1759_),
    .A2(_3473_),
    .Z(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7045_ (.A1(_2729_),
    .A2(_2874_),
    .Z(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7046_ (.A1(_0328_),
    .A2(_3459_),
    .A3(_2812_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7047_ (.A1(_2875_),
    .A2(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _7048_ (.A1(_2868_),
    .A2(_2873_),
    .A3(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _7049_ (.A1(_2859_),
    .A2(_2863_),
    .A3(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7050_ (.A1(_2858_),
    .A2(_2879_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7051_ (.A1(_2793_),
    .A2(_2797_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7052_ (.A1(_2798_),
    .A2(_2818_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7053_ (.A1(_2881_),
    .A2(_2882_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7054_ (.A1(_2880_),
    .A2(_2883_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7055_ (.I(_2833_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7056_ (.A1(_2885_),
    .A2(_2834_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7057_ (.A1(_2835_),
    .A2(_2836_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7058_ (.A1(_2886_),
    .A2(_2887_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7059_ (.A1(_2803_),
    .A2(_2816_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7060_ (.A1(_2802_),
    .A2(_2817_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7061_ (.A1(_2889_),
    .A2(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7062_ (.A1(_0343_),
    .A2(_3451_),
    .A3(_2724_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7063_ (.I(_1634_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7064_ (.A1(_2893_),
    .A2(_3434_),
    .A3(_2807_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7065_ (.A1(_2892_),
    .A2(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7066_ (.A1(_0354_),
    .A2(_3435_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7067_ (.A1(_2895_),
    .A2(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7068_ (.A1(_1519_),
    .A2(_3427_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7069_ (.A1(_2897_),
    .A2(_2898_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7070_ (.A1(_2891_),
    .A2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7071_ (.A1(_2888_),
    .A2(_2900_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7072_ (.A1(_2884_),
    .A2(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7073_ (.I(_2819_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7074_ (.A1(_2903_),
    .A2(_2822_),
    .Z(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7075_ (.A1(_2823_),
    .A2(_2839_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7076_ (.A1(_2904_),
    .A2(_2905_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7077_ (.A1(_2902_),
    .A2(_2906_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7078_ (.A1(_2830_),
    .A2(_2837_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7079_ (.A1(_2827_),
    .A2(_2838_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7080_ (.A1(_2908_),
    .A2(_2909_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7081_ (.I(_2910_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7082_ (.A1(_2907_),
    .A2(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7083_ (.A1(_2840_),
    .A2(_2843_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7084_ (.A1(_2840_),
    .A2(_2843_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7085_ (.A1(_2914_),
    .A2(_2846_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7086_ (.A1(_2913_),
    .A2(_2915_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7087_ (.A1(_2912_),
    .A2(_2916_),
    .Z(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7088_ (.A1(_2912_),
    .A2(_2916_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7089_ (.I(_2918_),
    .Z(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7090_ (.A1(_2917_),
    .A2(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _7091_ (.A1(_2239_),
    .A2(_2348_),
    .A3(_2441_),
    .A4(_2542_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _7092_ (.A1(_2616_),
    .A2(_2698_),
    .A3(_2771_),
    .A4(_2850_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7093_ (.A1(_2921_),
    .A2(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7094_ (.A1(_2774_),
    .A2(_2776_),
    .B(_2850_),
    .C(_2771_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7095_ (.A1(_2786_),
    .A2(_2848_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7096_ (.A1(_2849_),
    .A2(_2924_),
    .A3(_2925_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7097_ (.A1(_2619_),
    .A2(_2622_),
    .B(_2922_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7098_ (.A1(_2923_),
    .A2(_2926_),
    .A3(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _7099_ (.A1(_2242_),
    .A2(_2245_),
    .A3(_2926_),
    .A4(_2927_),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7100_ (.A1(_2250_),
    .A2(_2929_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7101_ (.A1(_2928_),
    .A2(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7102_ (.A1(_2920_),
    .A2(_2931_),
    .Z(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7103_ (.I0(\dspArea_regP[32] ),
    .I1(_2932_),
    .S(_2628_),
    .Z(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7104_ (.A1(_2856_),
    .A2(_2933_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7105_ (.I(\dspArea_regP[33] ),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7106_ (.A1(_2920_),
    .A2(_2931_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7107_ (.A1(_2902_),
    .A2(_2906_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7108_ (.A1(_2907_),
    .A2(_2911_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7109_ (.A1(_2936_),
    .A2(_2937_),
    .Z(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7110_ (.A1(_1759_),
    .A2(_3479_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7111_ (.A1(_1333_),
    .A2(_3473_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7112_ (.A1(_2939_),
    .A2(_2940_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7113_ (.A1(_2874_),
    .A2(_2870_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7114_ (.A1(_2871_),
    .A2(_2872_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7115_ (.A1(_2942_),
    .A2(_2943_),
    .Z(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7116_ (.A1(_2941_),
    .A2(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7117_ (.A1(_1634_),
    .A2(_3451_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7118_ (.A1(_0915_),
    .A2(_3458_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7119_ (.A1(_0333_),
    .A2(_3466_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7120_ (.A1(_2947_),
    .A2(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7121_ (.A1(_2946_),
    .A2(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7122_ (.A1(_2945_),
    .A2(_2950_),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7123_ (.A1(_2875_),
    .A2(_2876_),
    .B(_2873_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7124_ (.A1(_2875_),
    .A2(_2876_),
    .A3(_2873_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7125_ (.A1(_2868_),
    .A2(_2953_),
    .A3(_2952_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7126_ (.A1(_2952_),
    .A2(_2954_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7127_ (.A1(_2951_),
    .A2(_2955_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7128_ (.A1(_2934_),
    .A2(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7129_ (.A1(\dspArea_regP[32] ),
    .A2(_2857_),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7130_ (.A1(_2858_),
    .A2(_2879_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7131_ (.A1(_2958_),
    .A2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7132_ (.A1(_2957_),
    .A2(_2960_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7133_ (.I(_2895_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7134_ (.A1(_2962_),
    .A2(_2896_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7135_ (.A1(_2897_),
    .A2(_2898_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7136_ (.A1(_2963_),
    .A2(_2964_),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7137_ (.A1(_2860_),
    .A2(_2861_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7138_ (.A1(_2862_),
    .A2(_2966_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7139_ (.A1(_2859_),
    .A2(_2878_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7140_ (.A1(_2859_),
    .A2(_2878_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7141_ (.A1(_2967_),
    .A2(_2968_),
    .B(_2969_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7142_ (.A1(_1414_),
    .A2(_3459_),
    .A3(_2806_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7143_ (.A1(_1416_),
    .A2(_3443_),
    .A3(_2867_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7144_ (.A1(_2971_),
    .A2(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7145_ (.A1(_1847_),
    .A2(_3444_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7146_ (.A1(_2973_),
    .A2(_2974_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7147_ (.A1(_1297_),
    .A2(_3435_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7148_ (.A1(_2975_),
    .A2(_2976_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7149_ (.A1(_2970_),
    .A2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7150_ (.A1(_2965_),
    .A2(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7151_ (.A1(_2961_),
    .A2(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7152_ (.I(_2880_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7153_ (.A1(_2981_),
    .A2(_2883_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7154_ (.A1(_2884_),
    .A2(_2901_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7155_ (.A1(_2982_),
    .A2(_2983_),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7156_ (.A1(_2980_),
    .A2(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7157_ (.A1(_2891_),
    .A2(_2899_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7158_ (.A1(_2888_),
    .A2(_2900_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7159_ (.A1(_2986_),
    .A2(_2987_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7160_ (.A1(_2985_),
    .A2(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7161_ (.A1(_2938_),
    .A2(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7162_ (.A1(_2919_),
    .A2(_2935_),
    .A3(_2990_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7163_ (.A1(_2919_),
    .A2(_2935_),
    .B(_2990_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7164_ (.A1(_1831_),
    .A2(_2991_),
    .A3(_2992_),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7165_ (.A1(_2934_),
    .A2(_2454_),
    .B(_2993_),
    .C(_2855_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7166_ (.A1(\dspArea_regP[33] ),
    .A2(_2956_),
    .Z(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7167_ (.A1(_1845_),
    .A2(_3460_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7168_ (.A1(_0342_),
    .A2(_3467_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7169_ (.A1(_0334_),
    .A2(_3474_),
    .Z(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7170_ (.A1(_2996_),
    .A2(_2997_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7171_ (.A1(_2995_),
    .A2(_2998_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7172_ (.A1(_0328_),
    .A2(_3481_),
    .A3(_2869_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7173_ (.A1(_2999_),
    .A2(_3000_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7174_ (.I(_2944_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7175_ (.A1(_2941_),
    .A2(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7176_ (.A1(_2945_),
    .A2(_2950_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7177_ (.A1(_3003_),
    .A2(_3004_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7178_ (.A1(_3001_),
    .A2(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7179_ (.A1(\dspArea_regP[34] ),
    .A2(_3006_),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7180_ (.A1(_2994_),
    .A2(_3007_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7181_ (.I(_2973_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7182_ (.A1(_3009_),
    .A2(_2974_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7183_ (.A1(_2975_),
    .A2(_2976_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7184_ (.A1(_3010_),
    .A2(_3011_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7185_ (.I(_2951_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7186_ (.A1(_3013_),
    .A2(_2955_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7187_ (.A1(_0343_),
    .A2(_3468_),
    .A3(_2866_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7188_ (.A1(_1845_),
    .A2(_3451_),
    .A3(_2949_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7189_ (.A1(_3015_),
    .A2(_3016_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7190_ (.A1(_1847_),
    .A2(_3452_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7191_ (.A1(_3017_),
    .A2(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7192_ (.A1(_1519_),
    .A2(_3444_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7193_ (.A1(_3019_),
    .A2(_3020_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7194_ (.A1(_3014_),
    .A2(_3021_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7195_ (.A1(_3012_),
    .A2(_3022_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7196_ (.A1(_3008_),
    .A2(_3023_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7197_ (.I(_2960_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7198_ (.A1(_2957_),
    .A2(_3025_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7199_ (.A1(_2961_),
    .A2(_2979_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7200_ (.A1(_3026_),
    .A2(_3027_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7201_ (.A1(_3024_),
    .A2(_3028_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7202_ (.A1(_2970_),
    .A2(_2977_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7203_ (.A1(_2965_),
    .A2(_2978_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7204_ (.A1(_3030_),
    .A2(_3031_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7205_ (.A1(_3029_),
    .A2(_3032_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7206_ (.A1(_2980_),
    .A2(_2984_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7207_ (.A1(_2985_),
    .A2(_2988_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7208_ (.A1(_3034_),
    .A2(_3035_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7209_ (.A1(_3033_),
    .A2(_3036_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7210_ (.A1(_2938_),
    .A2(_2989_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7211_ (.A1(_2938_),
    .A2(_2989_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7212_ (.A1(_2919_),
    .A2(_3039_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7213_ (.A1(_2917_),
    .A2(_2918_),
    .A3(_2990_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7214_ (.I(_3041_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7215_ (.A1(_2249_),
    .A2(_2929_),
    .B(_3042_),
    .C(_2928_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7216_ (.A1(_3038_),
    .A2(_3040_),
    .A3(_3043_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7217_ (.A1(_3037_),
    .A2(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7218_ (.I0(\dspArea_regP[34] ),
    .I1(_3045_),
    .S(_2628_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7219_ (.A1(_2856_),
    .A2(_3046_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7220_ (.I(\dspArea_regP[35] ),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7221_ (.A1(_3024_),
    .A2(_3028_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7222_ (.A1(_3029_),
    .A2(_3032_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7223_ (.A1(\dspArea_regP[34] ),
    .A2(_3006_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7224_ (.A1(_0350_),
    .A2(_3469_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7225_ (.A1(_1413_),
    .A2(_3474_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7226_ (.A1(_0334_),
    .A2(_3480_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7227_ (.A1(_3052_),
    .A2(_3053_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7228_ (.A1(_3051_),
    .A2(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7229_ (.A1(_2874_),
    .A2(_2999_),
    .B(_0328_),
    .C(_3482_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7230_ (.A1(_3055_),
    .A2(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7231_ (.A1(_3047_),
    .A2(_3057_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7232_ (.A1(_3050_),
    .A2(_3058_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7233_ (.I(_3017_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7234_ (.A1(_3060_),
    .A2(_3018_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7235_ (.A1(_3019_),
    .A2(_3020_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7236_ (.A1(_3061_),
    .A2(_3062_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7237_ (.I(_3001_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7238_ (.A1(_3064_),
    .A2(_3005_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7239_ (.A1(_2948_),
    .A2(_3052_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7240_ (.A1(_2893_),
    .A2(_3460_),
    .A3(_2998_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7241_ (.A1(_0354_),
    .A2(_3460_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7242_ (.A1(_3066_),
    .A2(_3067_),
    .A3(_3068_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7243_ (.A1(_3066_),
    .A2(_3067_),
    .B(_3068_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7244_ (.A1(_3069_),
    .A2(_3070_),
    .Z(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7245_ (.A1(_0360_),
    .A2(_3452_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7246_ (.A1(_3071_),
    .A2(_3072_),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7247_ (.A1(_3065_),
    .A2(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7248_ (.A1(_3063_),
    .A2(_3074_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7249_ (.A1(_3059_),
    .A2(_3075_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7250_ (.A1(_2994_),
    .A2(_3007_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7251_ (.A1(_3008_),
    .A2(_3023_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7252_ (.A1(_3077_),
    .A2(_3078_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7253_ (.A1(_3014_),
    .A2(_3021_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7254_ (.A1(_3012_),
    .A2(_3022_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7255_ (.A1(_3080_),
    .A2(_3081_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _7256_ (.A1(_3076_),
    .A2(_3079_),
    .A3(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7257_ (.A1(_3048_),
    .A2(_3049_),
    .A3(_3083_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7258_ (.A1(_3048_),
    .A2(_3049_),
    .B(_3083_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7259_ (.A1(_3084_),
    .A2(_3085_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7260_ (.I(_3037_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7261_ (.A1(_3033_),
    .A2(_3036_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7262_ (.A1(_3087_),
    .A2(_3044_),
    .B(_3088_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7263_ (.A1(_3086_),
    .A2(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7264_ (.A1(_0988_),
    .A2(_3090_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7265_ (.A1(_3047_),
    .A2(_2454_),
    .B(_3091_),
    .C(_2855_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7266_ (.A1(_3037_),
    .A2(_3041_),
    .A3(_3086_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7267_ (.A1(_2249_),
    .A2(_2929_),
    .B(_3092_),
    .C(_2928_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7268_ (.A1(_2918_),
    .A2(_3038_),
    .B(_3039_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7269_ (.A1(_3037_),
    .A2(_3086_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7270_ (.I(_3084_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7271_ (.A1(_3088_),
    .A2(_3096_),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _7272_ (.A1(_3094_),
    .A2(_3095_),
    .B(_3097_),
    .C(_3085_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7273_ (.A1(\dspArea_regP[35] ),
    .A2(_3057_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7274_ (.A1(_0343_),
    .A2(_3482_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7275_ (.A1(_0350_),
    .A2(_3474_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7276_ (.A1(_3100_),
    .A2(_3101_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7277_ (.A1(\dspArea_regP[36] ),
    .A2(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7278_ (.A1(_3099_),
    .A2(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7279_ (.A1(_3071_),
    .A2(_3072_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7280_ (.A1(_3070_),
    .A2(_3105_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7281_ (.I(_3056_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7282_ (.A1(_3055_),
    .A2(_3107_),
    .Z(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7283_ (.A1(_0335_),
    .A2(_3481_),
    .A3(_3052_),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7284_ (.A1(_2893_),
    .A2(_3468_),
    .A3(_3054_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7285_ (.A1(_0354_),
    .A2(_3468_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7286_ (.A1(_3109_),
    .A2(_3110_),
    .A3(_3111_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7287_ (.A1(_3109_),
    .A2(_3110_),
    .B(_3111_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7288_ (.A1(_3112_),
    .A2(_3113_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7289_ (.A1(_0360_),
    .A2(_3461_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7290_ (.A1(_3114_),
    .A2(_3115_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7291_ (.A1(_3108_),
    .A2(_3116_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7292_ (.A1(_3106_),
    .A2(_3117_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7293_ (.A1(_3104_),
    .A2(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7294_ (.A1(_3050_),
    .A2(_3058_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7295_ (.A1(_3059_),
    .A2(_3075_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7296_ (.A1(_3120_),
    .A2(_3121_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7297_ (.A1(_3119_),
    .A2(_3122_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7298_ (.A1(_3065_),
    .A2(_3073_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7299_ (.A1(_3063_),
    .A2(_3074_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7300_ (.A1(_3124_),
    .A2(_3125_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7301_ (.A1(_3123_),
    .A2(_3126_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7302_ (.A1(_3076_),
    .A2(_3079_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7303_ (.A1(_3076_),
    .A2(_3079_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7304_ (.A1(_3129_),
    .A2(_3082_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7305_ (.A1(_3128_),
    .A2(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7306_ (.A1(_3127_),
    .A2(_3131_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7307_ (.A1(_3093_),
    .A2(_3098_),
    .B(_3132_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7308_ (.A1(_3132_),
    .A2(_3093_),
    .A3(_3098_),
    .Z(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7309_ (.A1(_3133_),
    .A2(_3134_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7310_ (.A1(\dspArea_regP[36] ),
    .A2(_0380_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7311_ (.A1(_0451_),
    .A2(_3135_),
    .B(_3136_),
    .C(_2855_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7312_ (.A1(\dspArea_regP[37] ),
    .A2(_1085_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7313_ (.I(_3127_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7314_ (.A1(_3138_),
    .A2(_3131_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7315_ (.A1(_3139_),
    .A2(_3133_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7316_ (.I(_3122_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7317_ (.A1(_3119_),
    .A2(_3141_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7318_ (.A1(_3123_),
    .A2(_3126_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7319_ (.A1(\dspArea_regP[36] ),
    .A2(_3102_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7320_ (.A1(_2893_),
    .A2(_3482_),
    .Z(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7321_ (.A1(\dspArea_regP[37] ),
    .A2(_3145_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7322_ (.A1(_3144_),
    .A2(_3146_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7323_ (.A1(_0355_),
    .A2(_3475_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7324_ (.A1(_3052_),
    .A2(_3145_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7325_ (.I0(_3148_),
    .I1(_0355_),
    .S(_3149_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7326_ (.A1(_1406_),
    .A2(_3469_),
    .Z(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7327_ (.A1(_3150_),
    .A2(_3151_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7328_ (.A1(_0362_),
    .A2(_3461_),
    .A3(_3114_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7329_ (.A1(_3113_),
    .A2(_3153_),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7330_ (.A1(_3152_),
    .A2(_3154_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7331_ (.A1(_3147_),
    .A2(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7332_ (.A1(_3099_),
    .A2(_3103_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7333_ (.I(_3104_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7334_ (.A1(_3158_),
    .A2(_3118_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7335_ (.A1(_3157_),
    .A2(_3159_),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7336_ (.A1(_3156_),
    .A2(_3160_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7337_ (.A1(_3108_),
    .A2(_3116_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7338_ (.I(_3106_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7339_ (.A1(_3163_),
    .A2(_3117_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7340_ (.A1(_3162_),
    .A2(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7341_ (.A1(_3161_),
    .A2(_3165_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7342_ (.A1(_3142_),
    .A2(_3143_),
    .A3(_3166_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7343_ (.A1(_3142_),
    .A2(_3143_),
    .B(_3166_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7344_ (.A1(_3167_),
    .A2(_3168_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7345_ (.A1(_3140_),
    .A2(_3169_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7346_ (.A1(_0799_),
    .A2(_3170_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7347_ (.A1(_3498_),
    .A2(_3137_),
    .A3(_3171_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7348_ (.I(_3154_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7349_ (.A1(_3152_),
    .A2(_3172_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7350_ (.A1(\dspArea_regP[37] ),
    .A2(_3145_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7351_ (.A1(\dspArea_regP[38] ),
    .A2(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7352_ (.A1(_0356_),
    .A2(_3483_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7353_ (.A1(_0360_),
    .A2(_3475_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7354_ (.A1(_3176_),
    .A2(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7355_ (.A1(_0356_),
    .A2(_3149_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7356_ (.I(_3150_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7357_ (.A1(_3180_),
    .A2(_3151_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7358_ (.A1(_3179_),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7359_ (.A1(_3178_),
    .A2(_3182_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7360_ (.A1(_3175_),
    .A2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7361_ (.A1(_3144_),
    .A2(_3146_),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7362_ (.A1(_3147_),
    .A2(_3155_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7363_ (.A1(_3185_),
    .A2(_3186_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7364_ (.A1(_3184_),
    .A2(_3187_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7365_ (.A1(_3173_),
    .A2(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7366_ (.A1(_3156_),
    .A2(_3160_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7367_ (.A1(_3161_),
    .A2(_3165_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7368_ (.A1(_3190_),
    .A2(_3191_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7369_ (.A1(_3189_),
    .A2(_3192_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7370_ (.A1(_3139_),
    .A2(_3168_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7371_ (.A1(_3133_),
    .A2(_3194_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7372_ (.A1(_3167_),
    .A2(_3195_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7373_ (.A1(_3193_),
    .A2(_3196_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7374_ (.A1(\dspArea_regP[38] ),
    .A2(_0426_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7375_ (.A1(_0495_),
    .A2(_3197_),
    .B(_3198_),
    .C(_3521_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7376_ (.I(\dspArea_regP[39] ),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7377_ (.A1(_3189_),
    .A2(_3192_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7378_ (.I(_3167_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7379_ (.A1(_3133_),
    .A2(_3194_),
    .B(_3193_),
    .C(_3201_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7380_ (.A1(_3178_),
    .A2(_3182_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7381_ (.A1(_0362_),
    .A2(_3483_),
    .A3(_3148_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7382_ (.A1(\dspArea_regP[39] ),
    .A2(_3204_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7383_ (.A1(\dspArea_regP[38] ),
    .A2(_3174_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7384_ (.A1(_3175_),
    .A2(_3183_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7385_ (.A1(_3206_),
    .A2(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7386_ (.A1(_3205_),
    .A2(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7387_ (.A1(_3203_),
    .A2(_3209_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7388_ (.A1(_3173_),
    .A2(_3188_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7389_ (.A1(_3184_),
    .A2(_3187_),
    .B(_3211_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7390_ (.A1(_3210_),
    .A2(_3212_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7391_ (.A1(_3210_),
    .A2(_3212_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7392_ (.A1(_3213_),
    .A2(_3214_),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7393_ (.A1(_3200_),
    .A2(_3202_),
    .B(_3215_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _7394_ (.A1(_3200_),
    .A2(_3202_),
    .A3(_3215_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7395_ (.A1(_0379_),
    .A2(_3216_),
    .A3(_3217_),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7396_ (.A1(_3199_),
    .A2(_0423_),
    .B(_3218_),
    .C(_3521_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7397_ (.A1(_3193_),
    .A2(_3215_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7398_ (.A1(_3132_),
    .A2(_3169_),
    .A3(_3219_),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7399_ (.A1(_3098_),
    .A2(_3220_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7400_ (.A1(_3167_),
    .A2(_3219_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7401_ (.A1(_3200_),
    .A2(_3214_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7402_ (.A1(_3194_),
    .A2(_3222_),
    .B1(_3223_),
    .B2(_3213_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7403_ (.A1(_3093_),
    .A2(_3220_),
    .B(_3221_),
    .C(_3224_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7404_ (.A1(_3205_),
    .A2(_3208_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7405_ (.A1(_3203_),
    .A2(_3209_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7406_ (.A1(_3226_),
    .A2(_3227_),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7407_ (.I(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7408_ (.I(_0362_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7409_ (.A1(_3199_),
    .A2(_3148_),
    .B(_2795_),
    .C(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7410_ (.A1(\dspArea_regP[40] ),
    .A2(_3231_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7411_ (.A1(_3229_),
    .A2(_3232_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7412_ (.A1(_3225_),
    .A2(_3233_),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7413_ (.I0(\dspArea_regP[40] ),
    .I1(_3234_),
    .S(_0379_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7414_ (.A1(_2856_),
    .A2(_3235_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7415_ (.A1(\dspArea_regP[40] ),
    .A2(_3231_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7416_ (.A1(\dspArea_regP[41] ),
    .A2(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7417_ (.A1(\dspArea_regP[41] ),
    .A2(_3236_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7418_ (.A1(_3237_),
    .A2(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7419_ (.A1(_3229_),
    .A2(_3232_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7420_ (.A1(_3225_),
    .A2(_3233_),
    .B(_3240_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7421_ (.A1(_3239_),
    .A2(_3241_),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7422_ (.A1(\dspArea_regP[41] ),
    .A2(_0380_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7423_ (.A1(_0988_),
    .A2(_3242_),
    .B(_3243_),
    .C(_3521_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _7424_ (.A1(_3233_),
    .A2(_3239_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7425_ (.A1(_3240_),
    .A2(_3237_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7426_ (.A1(_3238_),
    .A2(_3245_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7427_ (.A1(_3225_),
    .A2(_3244_),
    .B(_3246_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7428_ (.A1(_0426_),
    .A2(_3247_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7429_ (.A1(_3365_),
    .A2(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _7430_ (.A1(_3365_),
    .A2(_0370_),
    .A3(_3247_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7431_ (.A1(_0154_),
    .A2(_3249_),
    .A3(_3250_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7432_ (.A1(\dspArea_regP[43] ),
    .A2(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7433_ (.A1(_2856_),
    .A2(_3251_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7434_ (.A1(\dspArea_regP[43] ),
    .A2(\dspArea_regP[42] ),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7435_ (.I(_3252_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7436_ (.A1(\dspArea_regP[43] ),
    .A2(_3365_),
    .A3(_3238_),
    .A4(_3245_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7437_ (.A1(_3225_),
    .A2(_3244_),
    .A3(_3253_),
    .B(_3254_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7438_ (.A1(_0369_),
    .A2(_3255_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7439_ (.A1(\dspArea_regP[44] ),
    .A2(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7440_ (.A1(_3492_),
    .A2(_3257_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _7441_ (.A1(\dspArea_regP[44] ),
    .A2(_0425_),
    .A3(_3247_),
    .A4(_3252_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7442_ (.A1(\dspArea_regP[45] ),
    .A2(_3258_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7443_ (.A1(\dspArea_regP[45] ),
    .A2(\dspArea_regP[44] ),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _7444_ (.A1(_0425_),
    .A2(_3247_),
    .A3(_3252_),
    .A4(_3260_),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7445_ (.A1(_0154_),
    .A2(_3259_),
    .A3(_3261_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7446_ (.A1(\dspArea_regP[46] ),
    .A2(_3261_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _7447_ (.A1(\dspArea_regP[46] ),
    .A2(_0370_),
    .A3(_3255_),
    .A4(_3260_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7448_ (.A1(_0154_),
    .A2(_3262_),
    .A3(_3263_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7449_ (.A1(\dspArea_regP[47] ),
    .A2(_3263_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _7450_ (.A1(_3489_),
    .A2(_3264_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7451_ (.D(_0125_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(_zz_1_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7452_ (.D(_0126_),
    .CLK(net202),
    .Q(\dacArea_dac_cnt_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7453_ (.D(_0127_),
    .CLK(net202),
    .Q(\dacArea_dac_cnt_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7454_ (.D(_0128_),
    .CLK(net202),
    .Q(\dacArea_dac_cnt_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7455_ (.D(_0129_),
    .CLK(net202),
    .Q(\dacArea_dac_cnt_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7456_ (.D(_0130_),
    .CLK(net200),
    .Q(\dacArea_dac_cnt_0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7457_ (.D(_0131_),
    .CLK(net200),
    .Q(\dacArea_dac_cnt_0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7458_ (.D(_0132_),
    .CLK(net201),
    .Q(\dacArea_dac_cnt_0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7459_ (.D(_0133_),
    .CLK(net201),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7460_ (.D(_0134_),
    .CLK(net200),
    .Q(\dacArea_dac_cnt_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7461_ (.D(_0135_),
    .CLK(net200),
    .Q(\dacArea_dac_cnt_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7462_ (.D(_0136_),
    .CLK(net203),
    .Q(\dacArea_dac_cnt_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7463_ (.D(_0137_),
    .CLK(net201),
    .Q(\dacArea_dac_cnt_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7464_ (.D(_0138_),
    .CLK(net203),
    .Q(\dacArea_dac_cnt_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7465_ (.D(_0139_),
    .CLK(net206),
    .Q(\dacArea_dac_cnt_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7466_ (.D(_0140_),
    .CLK(net204),
    .Q(\dacArea_dac_cnt_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7467_ (.D(_0141_),
    .CLK(net204),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7468_ (.D(_0142_),
    .CLK(net203),
    .Q(\dacArea_dac_cnt_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7469_ (.D(_0143_),
    .CLK(net205),
    .Q(\dacArea_dac_cnt_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7470_ (.D(_0144_),
    .CLK(net205),
    .Q(\dacArea_dac_cnt_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7471_ (.D(_0145_),
    .CLK(net203),
    .Q(\dacArea_dac_cnt_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7472_ (.D(_0146_),
    .CLK(net205),
    .Q(\dacArea_dac_cnt_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7473_ (.D(_0147_),
    .CLK(net206),
    .Q(\dacArea_dac_cnt_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7474_ (.D(_0148_),
    .CLK(net206),
    .Q(\dacArea_dac_cnt_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7475_ (.D(_0149_),
    .CLK(net204),
    .Q(net145));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7476_ (.D(_0150_),
    .CLK(net205),
    .Q(\dacArea_dac_cnt_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7477_ (.D(_0151_),
    .CLK(net210),
    .Q(\dacArea_dac_cnt_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7478_ (.D(_0152_),
    .CLK(net207),
    .Q(\dacArea_dac_cnt_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7479_ (.D(_0153_),
    .CLK(net207),
    .Q(\dacArea_dac_cnt_3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7480_ (.D(_0000_),
    .CLK(net211),
    .Q(\dacArea_dac_cnt_3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7481_ (.D(_0001_),
    .CLK(net211),
    .Q(\dacArea_dac_cnt_3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7482_ (.D(_0002_),
    .CLK(net215),
    .Q(\dacArea_dac_cnt_3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7483_ (.D(_0003_),
    .CLK(net206),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7484_ (.D(_0004_),
    .CLK(net210),
    .Q(\dacArea_dac_cnt_4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7485_ (.D(_0005_),
    .CLK(net210),
    .Q(\dacArea_dac_cnt_4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7486_ (.D(_0006_),
    .CLK(net212),
    .Q(\dacArea_dac_cnt_4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7487_ (.D(_0007_),
    .CLK(net212),
    .Q(\dacArea_dac_cnt_4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7488_ (.D(_0008_),
    .CLK(net210),
    .Q(\dacArea_dac_cnt_4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7489_ (.D(_0009_),
    .CLK(net213),
    .Q(\dacArea_dac_cnt_4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7490_ (.D(_0010_),
    .CLK(net213),
    .Q(\dacArea_dac_cnt_4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7491_ (.D(_0011_),
    .CLK(net213),
    .Q(net147));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7492_ (.D(_0012_),
    .CLK(net211),
    .Q(\dacArea_dac_cnt_5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7493_ (.D(_0013_),
    .CLK(net212),
    .Q(\dacArea_dac_cnt_5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7494_ (.D(_0014_),
    .CLK(net212),
    .Q(\dacArea_dac_cnt_5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7495_ (.D(_0015_),
    .CLK(net216),
    .Q(\dacArea_dac_cnt_5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7496_ (.D(_0016_),
    .CLK(net213),
    .Q(\dacArea_dac_cnt_5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7497_ (.D(_0017_),
    .CLK(net217),
    .Q(\dacArea_dac_cnt_5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7498_ (.D(_0018_),
    .CLK(net217),
    .Q(\dacArea_dac_cnt_5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7499_ (.D(_0019_),
    .CLK(net214),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7500_ (.D(_0020_),
    .CLK(net214),
    .Q(\dacArea_dac_cnt_6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7501_ (.D(_0021_),
    .CLK(net216),
    .Q(\dacArea_dac_cnt_6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7502_ (.D(_0022_),
    .CLK(net216),
    .Q(\dacArea_dac_cnt_6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7503_ (.D(_0023_),
    .CLK(net216),
    .Q(\dacArea_dac_cnt_6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7504_ (.D(_0024_),
    .CLK(net219),
    .Q(\dacArea_dac_cnt_6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7505_ (.D(_0025_),
    .CLK(net219),
    .Q(\dacArea_dac_cnt_6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7506_ (.D(_0026_),
    .CLK(net219),
    .Q(\dacArea_dac_cnt_6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7507_ (.D(_0027_),
    .CLK(net217),
    .Q(net150));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7508_ (.D(_0028_),
    .CLK(net219),
    .Q(\dacArea_dac_cnt_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7509_ (.D(_0029_),
    .CLK(net218),
    .Q(\dacArea_dac_cnt_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7510_ (.D(_0030_),
    .CLK(net220),
    .Q(\dacArea_dac_cnt_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7511_ (.D(_0031_),
    .CLK(net220),
    .Q(\dacArea_dac_cnt_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7512_ (.D(_0032_),
    .CLK(net218),
    .Q(\dacArea_dac_cnt_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7513_ (.D(_0033_),
    .CLK(net220),
    .Q(\dacArea_dac_cnt_7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7514_ (.D(_0034_),
    .CLK(net221),
    .Q(\dacArea_dac_cnt_7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7515_ (.D(_0035_),
    .CLK(net217),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7516_ (.D(_0036_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7517_ (.D(_0037_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7518_ (.D(_0038_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7519_ (.D(_0039_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7520_ (.D(_0040_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7521_ (.D(_0041_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7522_ (.D(_0042_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7523_ (.D(_0043_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7524_ (.D(_0044_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7525_ (.D(_0045_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7526_ (.D(_0046_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7527_ (.D(_0047_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regA[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7528_ (.D(_0048_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7529_ (.D(_0049_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7530_ (.D(_0050_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7531_ (.D(_0051_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regA[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7532_ (.D(_0052_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7533_ (.D(_0053_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7534_ (.D(_0054_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7535_ (.D(_0055_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7536_ (.D(_0056_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7537_ (.D(_0057_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7538_ (.D(_0058_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7539_ (.D(_0059_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7540_ (.D(_0060_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7541_ (.D(_0061_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7542_ (.D(_0062_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7543_ (.D(_0063_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7544_ (.D(_0064_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7545_ (.D(_0065_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7546_ (.D(_0066_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7547_ (.D(_0067_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7548_ (.D(_0068_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7549_ (.D(_0069_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7550_ (.D(_0070_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7551_ (.D(_0071_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7552_ (.D(_0072_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7553_ (.D(_0073_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regB[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7554_ (.D(_0074_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7555_ (.D(_0075_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regB[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7556_ (.D(_0076_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regB[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7557_ (.D(_0077_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7558_ (.D(_0078_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7559_ (.D(_0079_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7560_ (.D(_0080_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7561_ (.D(_0081_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7562_ (.D(_0082_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7563_ (.D(_0083_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7564_ (.D(_0084_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7565_ (.D(_0085_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7566_ (.D(_0086_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7567_ (.D(_0087_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7568_ (.D(_0088_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7569_ (.D(_0089_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7570_ (.D(_0090_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _7571_ (.D(_0091_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7572_ (.D(_0092_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7573_ (.D(_0093_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7574_ (.D(_0094_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7575_ (.D(_0095_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _7576_ (.D(_0096_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7577_ (.D(_0097_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7578_ (.D(_0098_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7579_ (.D(_0099_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7580_ (.D(_0100_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7581_ (.D(_0101_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7582_ (.D(_0102_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7583_ (.D(_0103_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7584_ (.D(_0104_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7585_ (.D(_0105_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7586_ (.D(_0106_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7587_ (.D(_0107_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7588_ (.D(_0108_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7589_ (.D(_0109_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7590_ (.D(_0110_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7591_ (.D(_0111_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7592_ (.D(_0112_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7593_ (.D(_0113_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7594_ (.D(_0114_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7595_ (.D(_0115_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7596_ (.D(_0116_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regP[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7597_ (.D(_0117_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7598_ (.D(_0118_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7599_ (.D(_0119_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7600_ (.D(_0120_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7601_ (.D(_0121_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7602_ (.D(_0122_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7603_ (.D(_0123_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7604_ (.D(_0124_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[47] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_231 (.Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_232 (.Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_233 (.Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_234 (.Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_235 (.Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_236 (.Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_237 (.Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_238 (.Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_239 (.Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_240 (.Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_241 (.Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_242 (.Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_243 (.Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_244 (.Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_245 (.Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_246 (.Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_247 (.Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_248 (.Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_249 (.Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_250 (.Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_251 (.Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_252 (.Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_253 (.Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_254 (.Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_255 (.Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_256 (.Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_257 (.Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_258 (.Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_259 (.Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_260 (.Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_261 (.Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_262 (.Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_263 (.Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_264 (.Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_265 (.Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_266 (.Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_267 (.Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_230 (.Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7649_ (.I(net199),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7650_ (.I(net198),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7651_ (.I(net197),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7652_ (.I(net196),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7653_ (.I(net195),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7654_ (.I(net194),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7655_ (.I(net193),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7656_ (.I(net192),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7657_ (.I(net199),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7658_ (.I(net198),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7659_ (.I(net197),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7660_ (.I(net196),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7661_ (.I(net195),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7662_ (.I(net194),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7663_ (.I(net193),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7664_ (.I(net192),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7665_ (.I(net199),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7666_ (.I(net198),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7667_ (.I(net197),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7668_ (.I(net196),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7669_ (.I(net195),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7670_ (.I(net194),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7671_ (.I(net193),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7672_ (.I(net192),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input1 (.I(la_data_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(la_data_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(la_data_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(la_data_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(la_data_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(la_data_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(la_data_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input8 (.I(la_data_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(la_data_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(la_data_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(la_data_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input12 (.I(la_data_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(la_data_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(la_data_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(la_data_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(la_data_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(la_data_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input18 (.I(la_data_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(la_data_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(la_data_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(la_data_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(la_data_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(la_data_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(la_data_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(la_data_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(la_data_in[32]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input27 (.I(la_data_in[33]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(la_data_in[34]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(la_data_in[35]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input30 (.I(la_data_in[36]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input31 (.I(la_data_in[37]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input32 (.I(la_data_in[38]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(la_data_in[39]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(la_data_in[3]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input35 (.I(la_data_in[40]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input36 (.I(la_data_in[41]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input37 (.I(la_data_in[42]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input38 (.I(la_data_in[43]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(la_data_in[44]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(la_data_in[45]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(la_data_in[46]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(la_data_in[47]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input43 (.I(la_data_in[48]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(la_data_in[49]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input45 (.I(la_data_in[4]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(la_data_in[50]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(la_data_in[51]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(la_data_in[52]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(la_data_in[53]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input50 (.I(la_data_in[54]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input51 (.I(la_data_in[55]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input52 (.I(la_data_in[56]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(la_data_in[57]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input54 (.I(la_data_in[58]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input55 (.I(la_data_in[59]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input56 (.I(la_data_in[5]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input57 (.I(la_data_in[60]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input58 (.I(la_data_in[61]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input59 (.I(la_data_in[62]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input60 (.I(la_data_in[63]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input61 (.I(la_data_in[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input62 (.I(la_data_in[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input63 (.I(la_data_in[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input64 (.I(la_data_in[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(user_clock2),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input66 (.I(wb_ADR[0]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input67 (.I(wb_ADR[10]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input68 (.I(wb_ADR[11]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input69 (.I(wb_ADR[12]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input70 (.I(wb_ADR[13]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input71 (.I(wb_ADR[14]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input72 (.I(wb_ADR[15]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input73 (.I(wb_ADR[16]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input74 (.I(wb_ADR[17]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input75 (.I(wb_ADR[18]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input76 (.I(wb_ADR[19]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input77 (.I(wb_ADR[1]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input78 (.I(wb_ADR[20]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input79 (.I(wb_ADR[21]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input80 (.I(wb_ADR[22]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input81 (.I(wb_ADR[23]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input82 (.I(wb_ADR[24]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input83 (.I(wb_ADR[25]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input84 (.I(wb_ADR[26]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input85 (.I(wb_ADR[27]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input86 (.I(wb_ADR[28]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input87 (.I(wb_ADR[29]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input88 (.I(wb_ADR[2]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input89 (.I(wb_ADR[30]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input90 (.I(wb_ADR[31]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input91 (.I(wb_ADR[3]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input92 (.I(wb_ADR[4]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input93 (.I(wb_ADR[5]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input94 (.I(wb_ADR[6]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input95 (.I(wb_ADR[7]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input96 (.I(wb_ADR[8]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input97 (.I(wb_ADR[9]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input98 (.I(wb_CYC),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input99 (.I(wb_DAT_MOSI[0]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input100 (.I(wb_DAT_MOSI[10]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input101 (.I(wb_DAT_MOSI[11]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input102 (.I(wb_DAT_MOSI[12]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input103 (.I(wb_DAT_MOSI[13]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input104 (.I(wb_DAT_MOSI[14]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input105 (.I(wb_DAT_MOSI[15]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input106 (.I(wb_DAT_MOSI[16]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input107 (.I(wb_DAT_MOSI[17]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input108 (.I(wb_DAT_MOSI[18]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input109 (.I(wb_DAT_MOSI[19]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input110 (.I(wb_DAT_MOSI[1]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input111 (.I(wb_DAT_MOSI[20]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input112 (.I(wb_DAT_MOSI[21]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input113 (.I(wb_DAT_MOSI[22]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input114 (.I(wb_DAT_MOSI[23]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input115 (.I(wb_DAT_MOSI[24]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input116 (.I(wb_DAT_MOSI[2]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input117 (.I(wb_DAT_MOSI[3]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input118 (.I(wb_DAT_MOSI[4]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input119 (.I(wb_DAT_MOSI[5]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input120 (.I(wb_DAT_MOSI[6]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input121 (.I(wb_DAT_MOSI[7]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input122 (.I(wb_DAT_MOSI[8]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input123 (.I(wb_DAT_MOSI[9]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input124 (.I(wb_STB),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input125 (.I(wb_WE),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input126 (.I(wb_rst_i),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output127 (.I(net127),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output128 (.I(net128),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output129 (.I(net129),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output130 (.I(net130),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output131 (.I(net131),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output132 (.I(net132),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output133 (.I(net133),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output144 (.I(net144),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output145 (.I(net145),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output146 (.I(net146),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output147 (.I(net147),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output148 (.I(net148),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output149 (.I(net149),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output150 (.I(net150),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output151 (.I(net151),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output152 (.I(net152),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output153 (.I(net153),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output154 (.I(net154),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output155 (.I(net155),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output156 (.I(net156),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output157 (.I(net157),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output158 (.I(net158),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output159 (.I(net159),
    .Z(wb_ACK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output160 (.I(net160),
    .Z(wb_DAT_MISO[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output161 (.I(net161),
    .Z(wb_DAT_MISO[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output162 (.I(net162),
    .Z(wb_DAT_MISO[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output163 (.I(net163),
    .Z(wb_DAT_MISO[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output164 (.I(net164),
    .Z(wb_DAT_MISO[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output165 (.I(net165),
    .Z(wb_DAT_MISO[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output166 (.I(net166),
    .Z(wb_DAT_MISO[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output167 (.I(net167),
    .Z(wb_DAT_MISO[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output168 (.I(net168),
    .Z(wb_DAT_MISO[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output169 (.I(net169),
    .Z(wb_DAT_MISO[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output170 (.I(net170),
    .Z(wb_DAT_MISO[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output171 (.I(net171),
    .Z(wb_DAT_MISO[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output172 (.I(net172),
    .Z(wb_DAT_MISO[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output173 (.I(net173),
    .Z(wb_DAT_MISO[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output174 (.I(net174),
    .Z(wb_DAT_MISO[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output175 (.I(net175),
    .Z(wb_DAT_MISO[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output176 (.I(net176),
    .Z(wb_DAT_MISO[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output177 (.I(net177),
    .Z(wb_DAT_MISO[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output178 (.I(net178),
    .Z(wb_DAT_MISO[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output179 (.I(net179),
    .Z(wb_DAT_MISO[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output180 (.I(net180),
    .Z(wb_DAT_MISO[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output181 (.I(net181),
    .Z(wb_DAT_MISO[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output182 (.I(net182),
    .Z(wb_DAT_MISO[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output183 (.I(net183),
    .Z(wb_DAT_MISO[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output184 (.I(net184),
    .Z(wb_DAT_MISO[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output185 (.I(net185),
    .Z(wb_DAT_MISO[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output186 (.I(net186),
    .Z(wb_DAT_MISO[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output187 (.I(net187),
    .Z(wb_DAT_MISO[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output188 (.I(net188),
    .Z(wb_DAT_MISO[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output189 (.I(net189),
    .Z(wb_DAT_MISO[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output190 (.I(net190),
    .Z(wb_DAT_MISO[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output191 (.I(net191),
    .Z(wb_DAT_MISO[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout192 (.I(net151),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout193 (.I(net150),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout194 (.I(net148),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout195 (.I(net147),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout196 (.I(net146),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout197 (.I(net145),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout198 (.I(net144),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout199 (.I(net143),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout200 (.I(net201),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout201 (.I(net209),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout202 (.I(net209),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout203 (.I(net208),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout204 (.I(net208),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout205 (.I(net207),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout206 (.I(net207),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout207 (.I(net208),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout208 (.I(net209),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout209 (.I(net223),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout210 (.I(net211),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout211 (.I(net215),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout212 (.I(net214),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout213 (.I(net214),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net215),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout215 (.I(net222),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout216 (.I(net218),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout217 (.I(net218),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout218 (.I(net221),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout219 (.I(net220),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout220 (.I(net221),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout221 (.I(net222),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout222 (.I(net223),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout223 (.I(net65),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__D (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__D (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__D (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__D (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__D (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__D (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__D (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__I (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__I (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__I (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A4 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A3 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__I (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__I (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__I (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__I (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__I (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__I (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__C (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__C (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__C (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__C (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__B (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__C (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__C (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__C (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__C (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__I (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__I (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__I (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__I0 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__I (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__I (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__I (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__I (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__I (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I0 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__I (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__I (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__I (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I0 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__I (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__I (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I0 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__I (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__I (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__I0 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__I0 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__I (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I0 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__I (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__I (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__I (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I0 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__I0 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I0 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__I (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__B (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__I0 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__I0 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__I (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I0 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__S (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__S (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__S (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__S (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__I (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__I0 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__I1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__I0 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I0 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A4 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__I (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__S (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__S (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__S (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__S (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__S (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__S (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__I (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A3 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__B (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__B (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__I (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A3 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__I (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A3 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A3 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__I (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A3 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A3 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A3 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A4 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A3 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A3 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__S (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__S (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__S (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__S (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__I (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A3 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A3 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A3 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__I1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A3 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A3 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__I (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A4 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A3 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__C (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A3 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A3 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A3 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__I (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__I1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__C (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A3 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A3 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A3 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__B (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A3 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__C (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__C (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__C (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__C (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__I (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A3 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A3 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A3 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A3 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__B (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A3 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__I (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A3 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A3 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A3 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__B (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A3 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__I (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__I (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A3 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A3 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A3 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__B (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__I1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A3 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A3 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A3 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__I (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A3 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__B (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__I (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A3 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A3 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A3 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A3 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__B (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A3 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A3 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__B (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A3 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__B (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__C (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__B (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__C (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__S (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__S (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__S (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__S (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A3 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A3 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A3 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A3 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A3 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__B (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A3 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A3 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A3 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__B (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A3 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A3 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A3 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A3 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A3 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A3 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__B (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A3 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A3 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A3 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A3 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A3 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A3 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I1 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A3 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__I (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A3 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A3 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A3 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A3 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A3 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__B (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__I (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A3 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A2 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A3 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__I (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A3 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A3 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__B (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A3 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__I (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A3 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A2 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A3 (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__I1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A1 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__I (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A2 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A3 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A3 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A3 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A3 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__B (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A3 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A3 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A3 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__B (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A3 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A3 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__I (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A3 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A3 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A3 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__B (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A3 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A3 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A4 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__B1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__C (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A1 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A1 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__I1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__C (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__B (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__I (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A3 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A3 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A3 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A3 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__B (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A3 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A3 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__I (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__B (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__C (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__C (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__C (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__C (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A3 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A3 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__I (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A3 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A3 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A1 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A2 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A2 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A2 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A3 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__B (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A3 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__B (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__A3 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__C (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__B (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__I (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A3 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__A3 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A3 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A3 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__B (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A1 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A3 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A4 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__B (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__I (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A2 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A2 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A2 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A3 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__B (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A3 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A1 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A1 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A3 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__B (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A3 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__B (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A3 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A3 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A3 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A3 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__I (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__I1 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__S (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__S (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__S (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__S (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A3 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A3 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__I (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A1 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A2 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A2 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A3 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A3 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A1 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__B (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A3 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A3 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A2 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A3 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__I (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__B (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A2 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A1 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A3 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A3 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A2 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A3 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A2 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__I (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A4 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__B (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A3 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A3 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A1 (.I(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A2 (.I(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__A1 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A4 (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A3 (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__C (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__C (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A1 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__I1 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A1 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__I (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A2 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A2 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A2 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__I (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A2 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A2 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__I (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A1 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A1 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A1 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A1 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A1 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I1 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A3 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__B (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A3 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A3 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A1 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__B (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A3 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A2 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A3 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A3 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A3 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A3 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A1 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A4 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__B1 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__B1 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__B1 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__I (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A3 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__B2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__I (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__I (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__C1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__C1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__C1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__I (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__B2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__I (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__I (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__B2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__I (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__I (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__B1 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__I (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__I (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__I (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__B2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__I (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__I (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A2 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__I (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__I (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__I (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__B2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__I (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__I (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__I (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B2 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A2 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__I (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__B2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__I (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__I (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__I (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__I (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__B2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A4 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__I (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__I (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__I (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__B2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A2 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A1 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__I (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__I (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__I (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__I (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__B2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__I (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__B1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__B1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__I (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A2 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__I (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__B2 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__C1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__C1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__C1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__C1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__I (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__I (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__I (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__I (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__B2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A2 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__I (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__I (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A2 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__I (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A2 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A2 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__I (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__I (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__I (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__I (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A2 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__A2 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__I (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A2 (.I(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__I (.I(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__I (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__I (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A2 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A2 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A2 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A2 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__B2 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__C1 (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A2 (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A2 (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A2 (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__I (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A2 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__I (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__I (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A2 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A1 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A2 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A2 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A2 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__I (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__I (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A2 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A2 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__I (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A1 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__I (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__I (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A2 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A2 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__I (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A2 (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A2 (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__I (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A2 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__I (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__I (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A2 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A2 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A2 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A2 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__I (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__I (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__I (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__I (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A2 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A2 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__I (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A2 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A2 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A2 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A2 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A2 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A2 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__I (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__I (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A2 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A2 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A2 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A2 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A2 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A3 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__I (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__I (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__I (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A3 (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__C (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__C (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__C (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__I (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__I (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__I (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__I (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A1 (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__B (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A3 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A3 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(\dacArea_dac_cnt_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(\dacArea_dac_cnt_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(\dacArea_dac_cnt_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__I (.I(\dspArea_regA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__I (.I(\dspArea_regA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A2 (.I(\dspArea_regA[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(\dspArea_regA[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__I (.I(\dspArea_regA[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(\dspArea_regA[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(\dspArea_regA[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__I (.I(\dspArea_regA[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(\dspArea_regA[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(\dspArea_regA[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__I (.I(\dspArea_regA[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(\dspArea_regA[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__I (.I(\dspArea_regA[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__I (.I(\dspArea_regA[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__I (.I(\dspArea_regA[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A2 (.I(\dspArea_regA[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__I (.I(\dspArea_regA[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(\dspArea_regA[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__I (.I(\dspArea_regA[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(\dspArea_regA[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__I (.I(\dspArea_regA[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(\dspArea_regA[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(\dspArea_regA[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(\dspArea_regA[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__I (.I(\dspArea_regA[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A2 (.I(\dspArea_regA[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(\dspArea_regA[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(\dspArea_regA[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__I (.I(\dspArea_regA[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A2 (.I(\dspArea_regA[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(\dspArea_regA[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(\dspArea_regA[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(\dspArea_regA[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(\dspArea_regA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__I (.I(\dspArea_regA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__I (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__I (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__I (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A2 (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A2 (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__I (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A2 (.I(\dspArea_regA[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(\dspArea_regA[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(\dspArea_regA[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(\dspArea_regA[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__I (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(\dspArea_regA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(\dspArea_regA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__I (.I(\dspArea_regA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(\dspArea_regA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(\dspArea_regA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(\dspArea_regA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(\dspArea_regA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(\dspArea_regA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A2 (.I(\dspArea_regA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__I (.I(\dspArea_regA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(\dspArea_regA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A2 (.I(\dspArea_regA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(\dspArea_regA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__I (.I(\dspArea_regA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A2 (.I(\dspArea_regA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(\dspArea_regA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(\dspArea_regA[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(\dspArea_regA[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__I (.I(\dspArea_regA[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(\dspArea_regA[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(\dspArea_regA[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(\dspArea_regA[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__I (.I(\dspArea_regA[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(\dspArea_regB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__I (.I(\dspArea_regB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__I (.I(\dspArea_regB[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I (.I(\dspArea_regB[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(\dspArea_regB[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(\dspArea_regB[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(\dspArea_regB[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A1 (.I(\dspArea_regB[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(\dspArea_regB[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I (.I(\dspArea_regB[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__I (.I(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I (.I(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__I (.I(\dspArea_regB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__I (.I(\dspArea_regB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__I (.I(\dspArea_regB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(\dspArea_regB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(\dspArea_regB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(\dspArea_regB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__I (.I(\dspArea_regB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__I (.I(\dspArea_regB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(\dspArea_regB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(\dspArea_regB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I (.I(\dspArea_regB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(\dspArea_regB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(\dspArea_regB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(\dspArea_regB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I (.I(\dspArea_regB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I (.I(\dspArea_regB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__I (.I(\dspArea_regB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A1 (.I(\dspArea_regB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(\dspArea_regB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__I (.I(\dspArea_regB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(\dspArea_regB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I (.I(\dspArea_regB[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__I (.I(\dspArea_regB[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__I (.I(\dspArea_regB[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__I (.I(\dspArea_regB[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I (.I(\dspArea_regB[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__I (.I(\dspArea_regB[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__C2 (.I(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__I0 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__C2 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__C2 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__I0 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__C2 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__C2 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__C2 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__C2 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__I0 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I0 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I0 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A1 (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__I (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A1 (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__I0 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__I0 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__I (.I(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__I (.I(\dspArea_regP[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(\dspArea_regP[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A1 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__I0 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A1 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A1 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I0 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__C2 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I0 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A1 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__I (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A1 (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__I0 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A1 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A1 (.I(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__I (.I(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A1 (.I(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A1 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I0 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A1 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A1 (.I(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__I (.I(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A1 (.I(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A1 (.I(\dspArea_regP[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(\dspArea_regP[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(\dspArea_regP[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(\dspArea_regP[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__I0 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__C2 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A1 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__I0 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A1 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A2 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A1 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A1 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A1 (.I(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A1 (.I(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A1 (.I(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A1 (.I(\dspArea_regP[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A1 (.I(\dspArea_regP[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__C2 (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__C2 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I0 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__C2 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__I0 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__C2 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__C2 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I0 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A1 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__C2 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(la_data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(la_data_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(la_data_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(la_data_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(la_data_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(la_data_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(la_data_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(la_data_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(la_data_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(la_data_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(la_data_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(la_data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(la_data_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(la_data_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(la_data_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(la_data_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(la_data_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(la_data_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(la_data_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(la_data_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(la_data_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(la_data_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(la_data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(la_data_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(la_data_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(la_data_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(la_data_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(la_data_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(la_data_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(la_data_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(la_data_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(la_data_in[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(la_data_in[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(la_data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(la_data_in[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(la_data_in[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(la_data_in[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(la_data_in[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(la_data_in[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(la_data_in[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(la_data_in[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(la_data_in[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(la_data_in[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(la_data_in[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(la_data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(la_data_in[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(la_data_in[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(la_data_in[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(la_data_in[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(la_data_in[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(la_data_in[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(la_data_in[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(la_data_in[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(la_data_in[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(la_data_in[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(la_data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(la_data_in[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(la_data_in[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(la_data_in[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(la_data_in[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(la_data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(la_data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(la_data_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(la_data_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(user_clock2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(wb_ADR[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(wb_ADR[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(wb_ADR[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(wb_ADR[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(wb_ADR[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(wb_ADR[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(wb_ADR[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(wb_ADR[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(wb_ADR[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(wb_ADR[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(wb_ADR[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(wb_ADR[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(wb_ADR[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(wb_ADR[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(wb_ADR[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(wb_ADR[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(wb_ADR[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(wb_ADR[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(wb_ADR[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(wb_ADR[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(wb_ADR[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(wb_ADR[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(wb_ADR[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(wb_ADR[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(wb_ADR[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(wb_ADR[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(wb_ADR[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(wb_ADR[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(wb_ADR[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(wb_ADR[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(wb_ADR[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(wb_ADR[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(wb_CYC));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(wb_DAT_MOSI[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(wb_DAT_MOSI[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(wb_DAT_MOSI[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(wb_DAT_MOSI[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(wb_DAT_MOSI[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(wb_DAT_MOSI[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(wb_DAT_MOSI[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(wb_DAT_MOSI[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(wb_DAT_MOSI[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(wb_DAT_MOSI[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(wb_DAT_MOSI[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(wb_DAT_MOSI[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(wb_DAT_MOSI[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(wb_DAT_MOSI[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(wb_DAT_MOSI[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(wb_DAT_MOSI[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(wb_DAT_MOSI[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(wb_DAT_MOSI[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(wb_DAT_MOSI[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(wb_DAT_MOSI[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(wb_DAT_MOSI[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(wb_DAT_MOSI[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(wb_DAT_MOSI[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(wb_DAT_MOSI[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(wb_DAT_MOSI[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(wb_STB));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(wb_WE));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A2 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A3 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__I1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__I1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__I1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__I1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__I1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__I1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__I1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__I1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout199_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout198_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout197_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout193_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A3 (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__I (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__CLK (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout200_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__CLK (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout206_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout205_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout203_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout204_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout201_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__CLK (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout213_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__CLK (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout214_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__CLK (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout217_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout216_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout219_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout220_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout221_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout222_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout209_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net230;
 assign io_oeb[10] = net240;
 assign io_oeb[11] = net241;
 assign io_oeb[12] = net242;
 assign io_oeb[13] = net243;
 assign io_oeb[14] = net244;
 assign io_oeb[15] = net245;
 assign io_oeb[16] = net246;
 assign io_oeb[17] = net247;
 assign io_oeb[18] = net248;
 assign io_oeb[19] = net249;
 assign io_oeb[1] = net231;
 assign io_oeb[20] = net250;
 assign io_oeb[21] = net251;
 assign io_oeb[22] = net252;
 assign io_oeb[23] = net253;
 assign io_oeb[24] = net254;
 assign io_oeb[25] = net255;
 assign io_oeb[26] = net256;
 assign io_oeb[27] = net257;
 assign io_oeb[28] = net258;
 assign io_oeb[29] = net259;
 assign io_oeb[2] = net232;
 assign io_oeb[30] = net260;
 assign io_oeb[31] = net261;
 assign io_oeb[32] = net262;
 assign io_oeb[33] = net263;
 assign io_oeb[34] = net264;
 assign io_oeb[35] = net265;
 assign io_oeb[36] = net266;
 assign io_oeb[37] = net267;
 assign io_oeb[3] = net233;
 assign io_oeb[4] = net234;
 assign io_oeb[5] = net235;
 assign io_oeb[6] = net236;
 assign io_oeb[7] = net237;
 assign io_oeb[8] = net238;
 assign io_oeb[9] = net239;
 assign io_out[32] = net224;
 assign io_out[33] = net225;
 assign io_out[34] = net226;
 assign io_out[35] = net227;
 assign io_out[36] = net228;
 assign io_out[37] = net229;
endmodule

