// This is the unpowered netlist.
module DSP48 (user_clock2,
    wb_ACK,
    wb_CYC,
    wb_SEL,
    wb_STB,
    wb_WE,
    wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    wb_ADR,
    wb_DAT_MISO,
    wb_DAT_MOSI);
 input user_clock2;
 output wb_ACK;
 input wb_CYC;
 input wb_SEL;
 input wb_STB;
 input wb_WE;
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 input [31:0] wb_ADR;
 output [31:0] wb_DAT_MISO;
 input [31:0] wb_DAT_MOSI;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _zz_1_;
 wire \dacArea_dac_cnt_0[0] ;
 wire \dacArea_dac_cnt_0[1] ;
 wire \dacArea_dac_cnt_0[2] ;
 wire \dacArea_dac_cnt_0[3] ;
 wire \dacArea_dac_cnt_0[4] ;
 wire \dacArea_dac_cnt_0[5] ;
 wire \dacArea_dac_cnt_0[6] ;
 wire \dacArea_dac_cnt_1[0] ;
 wire \dacArea_dac_cnt_1[1] ;
 wire \dacArea_dac_cnt_1[2] ;
 wire \dacArea_dac_cnt_1[3] ;
 wire \dacArea_dac_cnt_1[4] ;
 wire \dacArea_dac_cnt_1[5] ;
 wire \dacArea_dac_cnt_1[6] ;
 wire \dacArea_dac_cnt_2[0] ;
 wire \dacArea_dac_cnt_2[1] ;
 wire \dacArea_dac_cnt_2[2] ;
 wire \dacArea_dac_cnt_2[3] ;
 wire \dacArea_dac_cnt_2[4] ;
 wire \dacArea_dac_cnt_2[5] ;
 wire \dacArea_dac_cnt_2[6] ;
 wire \dacArea_dac_cnt_3[0] ;
 wire \dacArea_dac_cnt_3[1] ;
 wire \dacArea_dac_cnt_3[2] ;
 wire \dacArea_dac_cnt_3[3] ;
 wire \dacArea_dac_cnt_3[4] ;
 wire \dacArea_dac_cnt_3[5] ;
 wire \dacArea_dac_cnt_3[6] ;
 wire \dacArea_dac_cnt_4[0] ;
 wire \dacArea_dac_cnt_4[1] ;
 wire \dacArea_dac_cnt_4[2] ;
 wire \dacArea_dac_cnt_4[3] ;
 wire \dacArea_dac_cnt_4[4] ;
 wire \dacArea_dac_cnt_4[5] ;
 wire \dacArea_dac_cnt_4[6] ;
 wire \dacArea_dac_cnt_5[0] ;
 wire \dacArea_dac_cnt_5[1] ;
 wire \dacArea_dac_cnt_5[2] ;
 wire \dacArea_dac_cnt_5[3] ;
 wire \dacArea_dac_cnt_5[4] ;
 wire \dacArea_dac_cnt_5[5] ;
 wire \dacArea_dac_cnt_5[6] ;
 wire \dacArea_dac_cnt_6[0] ;
 wire \dacArea_dac_cnt_6[1] ;
 wire \dacArea_dac_cnt_6[2] ;
 wire \dacArea_dac_cnt_6[3] ;
 wire \dacArea_dac_cnt_6[4] ;
 wire \dacArea_dac_cnt_6[5] ;
 wire \dacArea_dac_cnt_6[6] ;
 wire \dacArea_dac_cnt_7[0] ;
 wire \dacArea_dac_cnt_7[1] ;
 wire \dacArea_dac_cnt_7[2] ;
 wire \dacArea_dac_cnt_7[3] ;
 wire \dacArea_dac_cnt_7[4] ;
 wire \dacArea_dac_cnt_7[5] ;
 wire \dacArea_dac_cnt_7[6] ;
 wire \dspArea_regA[0] ;
 wire \dspArea_regA[10] ;
 wire \dspArea_regA[11] ;
 wire \dspArea_regA[12] ;
 wire \dspArea_regA[13] ;
 wire \dspArea_regA[14] ;
 wire \dspArea_regA[15] ;
 wire \dspArea_regA[16] ;
 wire \dspArea_regA[17] ;
 wire \dspArea_regA[18] ;
 wire \dspArea_regA[19] ;
 wire \dspArea_regA[1] ;
 wire \dspArea_regA[20] ;
 wire \dspArea_regA[21] ;
 wire \dspArea_regA[22] ;
 wire \dspArea_regA[23] ;
 wire \dspArea_regA[24] ;
 wire \dspArea_regA[2] ;
 wire \dspArea_regA[3] ;
 wire \dspArea_regA[4] ;
 wire \dspArea_regA[5] ;
 wire \dspArea_regA[6] ;
 wire \dspArea_regA[7] ;
 wire \dspArea_regA[8] ;
 wire \dspArea_regA[9] ;
 wire \dspArea_regB[0] ;
 wire \dspArea_regB[10] ;
 wire \dspArea_regB[11] ;
 wire \dspArea_regB[12] ;
 wire \dspArea_regB[13] ;
 wire \dspArea_regB[14] ;
 wire \dspArea_regB[15] ;
 wire \dspArea_regB[1] ;
 wire \dspArea_regB[2] ;
 wire \dspArea_regB[3] ;
 wire \dspArea_regB[4] ;
 wire \dspArea_regB[5] ;
 wire \dspArea_regB[6] ;
 wire \dspArea_regB[7] ;
 wire \dspArea_regB[8] ;
 wire \dspArea_regB[9] ;
 wire \dspArea_regP[0] ;
 wire \dspArea_regP[10] ;
 wire \dspArea_regP[11] ;
 wire \dspArea_regP[12] ;
 wire \dspArea_regP[13] ;
 wire \dspArea_regP[14] ;
 wire \dspArea_regP[15] ;
 wire \dspArea_regP[16] ;
 wire \dspArea_regP[17] ;
 wire \dspArea_regP[18] ;
 wire \dspArea_regP[19] ;
 wire \dspArea_regP[1] ;
 wire \dspArea_regP[20] ;
 wire \dspArea_regP[21] ;
 wire \dspArea_regP[22] ;
 wire \dspArea_regP[23] ;
 wire \dspArea_regP[24] ;
 wire \dspArea_regP[25] ;
 wire \dspArea_regP[26] ;
 wire \dspArea_regP[27] ;
 wire \dspArea_regP[28] ;
 wire \dspArea_regP[29] ;
 wire \dspArea_regP[2] ;
 wire \dspArea_regP[30] ;
 wire \dspArea_regP[31] ;
 wire \dspArea_regP[32] ;
 wire \dspArea_regP[33] ;
 wire \dspArea_regP[34] ;
 wire \dspArea_regP[35] ;
 wire \dspArea_regP[36] ;
 wire \dspArea_regP[37] ;
 wire \dspArea_regP[38] ;
 wire \dspArea_regP[39] ;
 wire \dspArea_regP[3] ;
 wire \dspArea_regP[40] ;
 wire \dspArea_regP[41] ;
 wire \dspArea_regP[42] ;
 wire \dspArea_regP[43] ;
 wire \dspArea_regP[44] ;
 wire \dspArea_regP[45] ;
 wire \dspArea_regP[46] ;
 wire \dspArea_regP[47] ;
 wire \dspArea_regP[4] ;
 wire \dspArea_regP[5] ;
 wire \dspArea_regP[6] ;
 wire \dspArea_regP[7] ;
 wire \dspArea_regP[8] ;
 wire \dspArea_regP[9] ;
 wire net199;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net200;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net201;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire clknet_0_wb_clk_i;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3392_ (.A1(net124),
    .A2(_zz_1_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3393_ (.I(_2976_),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3394_ (.A1(net83),
    .A2(net82),
    .A3(net85),
    .A4(net84),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3395_ (.A1(net79),
    .A2(net78),
    .A3(net81),
    .A4(net80),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3396_ (.A1(net74),
    .A2(net73),
    .A3(net76),
    .A4(net75),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3397_ (.A1(net87),
    .A2(net86),
    .A3(net90),
    .A4(net89),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _3398_ (.A1(_2978_),
    .A2(_2979_),
    .A3(_2980_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3399_ (.A1(_2977_),
    .A2(_2981_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3400_ (.A1(net70),
    .A2(net69),
    .A3(net72),
    .A4(net71),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3401_ (.A1(net97),
    .A2(net96),
    .A3(net68),
    .A4(net67),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3402_ (.A1(net77),
    .A2(net66),
    .A3(_2983_),
    .A4(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3403_ (.A1(_2982_),
    .A2(_2985_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3404_ (.I(net92),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3405_ (.A1(net93),
    .A2(net95),
    .A3(net94),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3406_ (.A1(_2987_),
    .A2(_2988_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3407_ (.A1(net88),
    .A2(_2989_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3408_ (.A1(net91),
    .A2(_2986_),
    .A3(_2990_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3409_ (.I(_2991_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3410_ (.I(net88),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3411_ (.I(net91),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3412_ (.A1(_2993_),
    .A2(_2994_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3413_ (.A1(_2982_),
    .A2(_2985_),
    .A3(_2995_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3414_ (.A1(net92),
    .A2(_2988_),
    .Z(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3415_ (.A1(_2996_),
    .A2(_2997_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3416_ (.I(_2998_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3417_ (.I(\dspArea_regA[0] ),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3418_ (.I(_3000_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3419_ (.I(_3001_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3420_ (.A1(_2993_),
    .A2(net91),
    .A3(_2986_),
    .A4(_2989_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3421_ (.I(_3003_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3422_ (.A1(\dspArea_regP[32] ),
    .A2(_2992_),
    .B1(_2999_),
    .B2(_3002_),
    .C1(_3004_),
    .C2(\dspArea_regP[0] ),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3423_ (.I(_3005_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3424_ (.I(_2998_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3425_ (.I(\dspArea_regA[1] ),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3426_ (.I(_3007_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3427_ (.I(_3008_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3428_ (.A1(\dspArea_regP[33] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3009_),
    .C1(_3004_),
    .C2(\dspArea_regP[1] ),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3429_ (.I(_3010_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3430_ (.I(\dspArea_regA[2] ),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3431_ (.I(_3011_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3432_ (.I(_3012_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3433_ (.A1(\dspArea_regP[34] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3013_),
    .C1(_3004_),
    .C2(\dspArea_regP[2] ),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3434_ (.I(_3014_),
    .ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3435_ (.I(\dspArea_regA[3] ),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3436_ (.I(_3015_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3437_ (.I(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3438_ (.A1(\dspArea_regP[35] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3017_),
    .C1(_3004_),
    .C2(\dspArea_regP[3] ),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3439_ (.I(_3018_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3440_ (.I(\dspArea_regA[4] ),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3441_ (.I(_3019_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3442_ (.I(_3020_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3443_ (.I(_3003_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3444_ (.A1(\dspArea_regP[36] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3021_),
    .C1(_3022_),
    .C2(\dspArea_regP[4] ),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3445_ (.I(_3023_),
    .ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3446_ (.I(\dspArea_regA[5] ),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3447_ (.I(_3024_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3448_ (.I(_3025_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3449_ (.A1(\dspArea_regP[37] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3026_),
    .C1(_3022_),
    .C2(\dspArea_regP[5] ),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3450_ (.I(_3027_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3451_ (.I(\dspArea_regA[6] ),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3452_ (.I(_3028_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3453_ (.I(_3029_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3454_ (.A1(\dspArea_regP[38] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3030_),
    .C1(_3022_),
    .C2(\dspArea_regP[6] ),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3455_ (.I(_3031_),
    .ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3456_ (.I(\dspArea_regA[7] ),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3457_ (.I(_3032_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3458_ (.I(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3459_ (.A1(\dspArea_regP[39] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3034_),
    .C1(_3022_),
    .C2(\dspArea_regP[7] ),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3460_ (.I(_3035_),
    .ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3461_ (.I(\dspArea_regA[8] ),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3462_ (.I(_3036_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3463_ (.I(_3037_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3464_ (.A1(\dspArea_regP[40] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3038_),
    .C1(_3022_),
    .C2(\dspArea_regP[8] ),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3465_ (.I(_3039_),
    .ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3466_ (.I(\dspArea_regA[9] ),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3467_ (.I(_3040_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3468_ (.I(_3041_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3469_ (.A1(\dspArea_regP[41] ),
    .A2(_2992_),
    .B1(_3006_),
    .B2(_3042_),
    .C1(_3022_),
    .C2(\dspArea_regP[9] ),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3470_ (.I(_3043_),
    .ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3471_ (.I(\dspArea_regA[10] ),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3472_ (.I(_3044_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3473_ (.I(_3045_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3474_ (.A1(\dspArea_regP[42] ),
    .A2(_2991_),
    .B1(_3006_),
    .B2(_3046_),
    .C1(_3022_),
    .C2(\dspArea_regP[10] ),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3475_ (.I(_3047_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3476_ (.I(\dspArea_regA[11] ),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3477_ (.I(_3048_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3478_ (.I(_3049_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3479_ (.A1(\dspArea_regP[43] ),
    .A2(_2991_),
    .B1(_2998_),
    .B2(_3050_),
    .C1(_3022_),
    .C2(\dspArea_regP[11] ),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3480_ (.I(_3051_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3481_ (.I(\dspArea_regA[12] ),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3482_ (.I(_3052_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3483_ (.I(_3053_),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3484_ (.A1(\dspArea_regP[44] ),
    .A2(_2991_),
    .B1(_2998_),
    .B2(_3054_),
    .C1(_3022_),
    .C2(\dspArea_regP[12] ),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3485_ (.I(_3055_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3486_ (.I(\dspArea_regA[13] ),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3487_ (.I(_3056_),
    .Z(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3488_ (.I(_3057_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3489_ (.A1(\dspArea_regP[45] ),
    .A2(_2991_),
    .B1(_2998_),
    .B2(_3058_),
    .C1(_3022_),
    .C2(\dspArea_regP[13] ),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3490_ (.I(_3059_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3491_ (.I(\dspArea_regA[14] ),
    .Z(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3492_ (.I(_3060_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3493_ (.I(_3061_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3494_ (.A1(\dspArea_regP[46] ),
    .A2(_2991_),
    .B1(_2998_),
    .B2(_3062_),
    .C1(_3003_),
    .C2(\dspArea_regP[14] ),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3495_ (.I(_3063_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3496_ (.I(\dspArea_regA[15] ),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3497_ (.I(_3064_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3498_ (.I(_3065_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3499_ (.A1(\dspArea_regP[47] ),
    .A2(_2991_),
    .B1(_2998_),
    .B2(_3066_),
    .C1(_3003_),
    .C2(\dspArea_regP[15] ),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3500_ (.I(_3067_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3501_ (.I(\dspArea_regA[16] ),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3502_ (.I(_3068_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3503_ (.I(_3069_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3504_ (.A1(_3070_),
    .A2(_2999_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3505_ (.I(_3003_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3506_ (.A1(\dspArea_regP[16] ),
    .A2(_3072_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3507_ (.A1(_3071_),
    .A2(_3073_),
    .ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3508_ (.I(\dspArea_regA[17] ),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3509_ (.I(_3074_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3510_ (.I(_3075_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3511_ (.A1(_3076_),
    .A2(_2999_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3512_ (.A1(\dspArea_regP[17] ),
    .A2(_3072_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3513_ (.A1(_3077_),
    .A2(_3078_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3514_ (.I(\dspArea_regA[18] ),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3515_ (.I(_3079_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3516_ (.I(_3080_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3517_ (.A1(_3081_),
    .A2(_2999_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3518_ (.A1(\dspArea_regP[18] ),
    .A2(_3072_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3519_ (.A1(_3082_),
    .A2(_3083_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3520_ (.I(\dspArea_regA[19] ),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3521_ (.I(_3084_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3522_ (.I(_3085_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3523_ (.A1(_3086_),
    .A2(_2999_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3524_ (.A1(\dspArea_regP[19] ),
    .A2(_3004_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3525_ (.A1(_3087_),
    .A2(_3088_),
    .ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3526_ (.I(\dspArea_regA[20] ),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3527_ (.I(_3089_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3528_ (.A1(_3090_),
    .A2(_2999_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3529_ (.A1(\dspArea_regP[20] ),
    .A2(_3004_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3530_ (.A1(_3091_),
    .A2(_3092_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3531_ (.I(\dspArea_regA[21] ),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3532_ (.I(_3093_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3533_ (.A1(_3094_),
    .A2(_2999_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3534_ (.A1(\dspArea_regP[21] ),
    .A2(_3004_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3535_ (.A1(_3095_),
    .A2(_3096_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3536_ (.I(\dspArea_regA[22] ),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3537_ (.I(_3097_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3538_ (.A1(_3098_),
    .A2(_2999_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3539_ (.A1(\dspArea_regP[22] ),
    .A2(_3004_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3540_ (.A1(_3099_),
    .A2(_3100_),
    .ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3541_ (.I(\dspArea_regA[23] ),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3542_ (.I(_3101_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3543_ (.A1(_3102_),
    .A2(_2999_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3544_ (.A1(\dspArea_regP[23] ),
    .A2(_3004_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3545_ (.A1(_3103_),
    .A2(_3104_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3546_ (.I(\dspArea_regA[24] ),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3547_ (.I(_3105_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3548_ (.A1(_3106_),
    .A2(_2999_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3549_ (.A1(\dspArea_regP[24] ),
    .A2(_3004_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3550_ (.A1(_3107_),
    .A2(_3108_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3551_ (.A1(\dspArea_regP[25] ),
    .A2(_3072_),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3552_ (.A1(\dspArea_regP[26] ),
    .A2(_3072_),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3553_ (.A1(\dspArea_regP[27] ),
    .A2(_3072_),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3554_ (.A1(\dspArea_regP[28] ),
    .A2(_3072_),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3555_ (.A1(\dspArea_regP[29] ),
    .A2(_3072_),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3556_ (.A1(\dspArea_regP[30] ),
    .A2(_3072_),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3557_ (.A1(\dspArea_regP[31] ),
    .A2(_3072_),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3558_ (.I(net126),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3559_ (.I(_3109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3560_ (.I(_3110_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3561_ (.A1(net124),
    .A2(net98),
    .A3(_3111_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3562_ (.I(_3109_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3563_ (.A1(\dacArea_dac_cnt_0[0] ),
    .A2(net1),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3564_ (.A1(\dacArea_dac_cnt_0[0] ),
    .A2(net1),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3565_ (.A1(_3112_),
    .A2(_3113_),
    .A3(_3114_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3566_ (.A1(\dacArea_dac_cnt_0[1] ),
    .A2(net12),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3567_ (.A1(_3114_),
    .A2(_3115_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3568_ (.A1(_3114_),
    .A2(_3115_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3569_ (.A1(_3111_),
    .A2(_3116_),
    .A3(_3117_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3570_ (.I(_3110_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3571_ (.A1(\dacArea_dac_cnt_0[1] ),
    .A2(net12),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3572_ (.A1(_3119_),
    .A2(_3117_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3573_ (.A1(\dacArea_dac_cnt_0[2] ),
    .A2(net23),
    .A3(_3120_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3574_ (.A1(_3118_),
    .A2(_3121_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3575_ (.A1(\dacArea_dac_cnt_0[2] ),
    .A2(net23),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3576_ (.A1(_3120_),
    .A2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3577_ (.A1(\dacArea_dac_cnt_0[2] ),
    .A2(net23),
    .B(_3123_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3578_ (.A1(\dacArea_dac_cnt_0[3] ),
    .A2(net34),
    .A3(_3124_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3579_ (.A1(_3118_),
    .A2(_3125_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3580_ (.A1(\dacArea_dac_cnt_0[3] ),
    .A2(net34),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3581_ (.A1(\dacArea_dac_cnt_0[3] ),
    .A2(net34),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3582_ (.A1(_3126_),
    .A2(_3124_),
    .B(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3583_ (.A1(\dacArea_dac_cnt_0[4] ),
    .A2(net45),
    .A3(_3128_),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3584_ (.A1(_3118_),
    .A2(_3129_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3585_ (.A1(\dacArea_dac_cnt_0[4] ),
    .A2(net45),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3586_ (.A1(\dacArea_dac_cnt_0[4] ),
    .A2(net45),
    .B(_3128_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3587_ (.A1(_3130_),
    .A2(_3131_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3588_ (.A1(\dacArea_dac_cnt_0[5] ),
    .A2(net56),
    .A3(_3132_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3589_ (.A1(_3118_),
    .A2(_3133_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3590_ (.A1(\dacArea_dac_cnt_0[5] ),
    .A2(net56),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3591_ (.A1(_3134_),
    .A2(_3132_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3592_ (.A1(\dacArea_dac_cnt_0[5] ),
    .A2(net56),
    .B(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3593_ (.A1(\dacArea_dac_cnt_0[6] ),
    .A2(net61),
    .A3(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3594_ (.A1(_3118_),
    .A2(_3137_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3595_ (.A1(\dacArea_dac_cnt_0[6] ),
    .A2(net61),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3596_ (.A1(\dacArea_dac_cnt_0[6] ),
    .A2(net61),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3597_ (.A1(_3138_),
    .A2(_3136_),
    .B(_3139_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3598_ (.A1(net143),
    .A2(net62),
    .A3(_3140_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3599_ (.A1(_3112_),
    .A2(_3141_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3600_ (.I(_3109_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3601_ (.A1(\dacArea_dac_cnt_1[0] ),
    .A2(net63),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3602_ (.A1(\dacArea_dac_cnt_1[0] ),
    .A2(net63),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3603_ (.A1(_3142_),
    .A2(_3143_),
    .A3(_3144_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3604_ (.A1(\dacArea_dac_cnt_1[1] ),
    .A2(net64),
    .Z(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3605_ (.A1(_3144_),
    .A2(_3145_),
    .Z(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3606_ (.A1(_3144_),
    .A2(_3145_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3607_ (.A1(_3111_),
    .A2(_3146_),
    .A3(_3147_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3608_ (.A1(\dacArea_dac_cnt_1[1] ),
    .A2(net64),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3609_ (.A1(_3148_),
    .A2(_3147_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3610_ (.A1(\dacArea_dac_cnt_1[2] ),
    .A2(net2),
    .A3(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3611_ (.A1(_3118_),
    .A2(_3150_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3612_ (.A1(\dacArea_dac_cnt_1[2] ),
    .A2(net2),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3613_ (.A1(_3149_),
    .A2(_3151_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3614_ (.A1(\dacArea_dac_cnt_1[2] ),
    .A2(net2),
    .B(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3615_ (.A1(\dacArea_dac_cnt_1[3] ),
    .A2(net3),
    .A3(_3153_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3616_ (.A1(_3118_),
    .A2(_3154_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3617_ (.A1(\dacArea_dac_cnt_1[3] ),
    .A2(net3),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3618_ (.A1(\dacArea_dac_cnt_1[3] ),
    .A2(net3),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3619_ (.A1(_3155_),
    .A2(_3153_),
    .B(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3620_ (.A1(\dacArea_dac_cnt_1[4] ),
    .A2(net4),
    .A3(_3157_),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3621_ (.A1(_3118_),
    .A2(_3158_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3622_ (.A1(\dacArea_dac_cnt_1[4] ),
    .A2(net4),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3623_ (.A1(\dacArea_dac_cnt_1[4] ),
    .A2(net4),
    .B(_3157_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3624_ (.A1(_3159_),
    .A2(_3160_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3625_ (.A1(\dacArea_dac_cnt_1[5] ),
    .A2(net5),
    .A3(_3161_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3626_ (.A1(_3118_),
    .A2(_3162_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3627_ (.A1(\dacArea_dac_cnt_1[5] ),
    .A2(net5),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3628_ (.A1(_3163_),
    .A2(_3161_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3629_ (.A1(\dacArea_dac_cnt_1[5] ),
    .A2(net5),
    .B(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3630_ (.A1(\dacArea_dac_cnt_1[6] ),
    .A2(net6),
    .A3(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3631_ (.A1(_3118_),
    .A2(_3166_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3632_ (.A1(\dacArea_dac_cnt_1[6] ),
    .A2(net6),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3633_ (.A1(\dacArea_dac_cnt_1[6] ),
    .A2(net6),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3634_ (.A1(_3167_),
    .A2(_3165_),
    .B(_3168_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3635_ (.A1(net144),
    .A2(net7),
    .A3(_3169_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3636_ (.A1(_3112_),
    .A2(_3170_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3637_ (.A1(\dacArea_dac_cnt_2[0] ),
    .A2(net8),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3638_ (.A1(\dacArea_dac_cnt_2[0] ),
    .A2(net8),
    .Z(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3639_ (.A1(_3142_),
    .A2(_3171_),
    .A3(_3172_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3640_ (.I(_3110_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3641_ (.A1(\dacArea_dac_cnt_2[1] ),
    .A2(net9),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3642_ (.A1(_3172_),
    .A2(_3174_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3643_ (.A1(_3172_),
    .A2(_3174_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3644_ (.A1(_3173_),
    .A2(_3175_),
    .A3(_3176_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3645_ (.I(_3110_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3646_ (.A1(\dacArea_dac_cnt_2[1] ),
    .A2(net9),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3647_ (.A1(_3178_),
    .A2(_3176_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3648_ (.A1(\dacArea_dac_cnt_2[2] ),
    .A2(net10),
    .A3(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3649_ (.A1(_3177_),
    .A2(_3180_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3650_ (.A1(\dacArea_dac_cnt_2[2] ),
    .A2(net10),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3651_ (.A1(_3179_),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3652_ (.A1(\dacArea_dac_cnt_2[2] ),
    .A2(net10),
    .B(_3182_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3653_ (.A1(\dacArea_dac_cnt_2[3] ),
    .A2(net11),
    .A3(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3654_ (.A1(_3177_),
    .A2(_3184_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3655_ (.A1(\dacArea_dac_cnt_2[3] ),
    .A2(net11),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3656_ (.A1(\dacArea_dac_cnt_2[3] ),
    .A2(net11),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3657_ (.A1(_3185_),
    .A2(_3183_),
    .B(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3658_ (.A1(\dacArea_dac_cnt_2[4] ),
    .A2(net13),
    .A3(_3187_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3659_ (.A1(_3177_),
    .A2(_3188_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3660_ (.A1(\dacArea_dac_cnt_2[4] ),
    .A2(net13),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3661_ (.A1(\dacArea_dac_cnt_2[4] ),
    .A2(net13),
    .B(_3187_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3662_ (.A1(_3189_),
    .A2(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3663_ (.A1(\dacArea_dac_cnt_2[5] ),
    .A2(net14),
    .A3(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3664_ (.A1(_3177_),
    .A2(_3192_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3665_ (.A1(\dacArea_dac_cnt_2[5] ),
    .A2(net14),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3666_ (.A1(_3193_),
    .A2(_3191_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3667_ (.A1(\dacArea_dac_cnt_2[5] ),
    .A2(net14),
    .B(_3194_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3668_ (.A1(\dacArea_dac_cnt_2[6] ),
    .A2(net15),
    .A3(_3195_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3669_ (.A1(_3177_),
    .A2(_3196_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3670_ (.A1(\dacArea_dac_cnt_2[6] ),
    .A2(net15),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3671_ (.A1(\dacArea_dac_cnt_2[6] ),
    .A2(net15),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3672_ (.A1(_3197_),
    .A2(_3195_),
    .B(_3198_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3673_ (.A1(net145),
    .A2(net16),
    .A3(_3199_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3674_ (.A1(_3112_),
    .A2(_3200_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3675_ (.A1(\dacArea_dac_cnt_3[0] ),
    .A2(net17),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3676_ (.A1(\dacArea_dac_cnt_3[0] ),
    .A2(net17),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3677_ (.A1(_3142_),
    .A2(_3201_),
    .A3(_3202_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3678_ (.A1(\dacArea_dac_cnt_3[1] ),
    .A2(net18),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3679_ (.A1(_3202_),
    .A2(_3203_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3680_ (.A1(_3202_),
    .A2(_3203_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3681_ (.A1(_3173_),
    .A2(_3204_),
    .A3(_3205_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3682_ (.A1(\dacArea_dac_cnt_3[1] ),
    .A2(net18),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3683_ (.A1(_3206_),
    .A2(_3205_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3684_ (.A1(\dacArea_dac_cnt_3[2] ),
    .A2(net19),
    .A3(_3207_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3685_ (.A1(_3177_),
    .A2(_3208_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3686_ (.A1(\dacArea_dac_cnt_3[2] ),
    .A2(net19),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3687_ (.A1(_3207_),
    .A2(_3209_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3688_ (.A1(\dacArea_dac_cnt_3[2] ),
    .A2(net19),
    .B(_3210_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3689_ (.A1(\dacArea_dac_cnt_3[3] ),
    .A2(net20),
    .A3(_3211_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3690_ (.A1(_3177_),
    .A2(_3212_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3691_ (.A1(\dacArea_dac_cnt_3[3] ),
    .A2(net20),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3692_ (.A1(\dacArea_dac_cnt_3[3] ),
    .A2(net20),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3693_ (.A1(_3213_),
    .A2(_3211_),
    .B(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3694_ (.A1(\dacArea_dac_cnt_3[4] ),
    .A2(net21),
    .A3(_3215_),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3695_ (.A1(_3177_),
    .A2(_3216_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3696_ (.A1(\dacArea_dac_cnt_3[4] ),
    .A2(net21),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3697_ (.A1(\dacArea_dac_cnt_3[4] ),
    .A2(net21),
    .B(_3215_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3698_ (.A1(_3217_),
    .A2(_3218_),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3699_ (.A1(\dacArea_dac_cnt_3[5] ),
    .A2(net22),
    .A3(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3700_ (.A1(_3177_),
    .A2(_3220_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3701_ (.A1(\dacArea_dac_cnt_3[5] ),
    .A2(net22),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3702_ (.A1(_3221_),
    .A2(_3219_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3703_ (.A1(\dacArea_dac_cnt_3[5] ),
    .A2(net22),
    .B(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3704_ (.A1(\dacArea_dac_cnt_3[6] ),
    .A2(net24),
    .A3(_3223_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3705_ (.A1(_3177_),
    .A2(_3224_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3706_ (.A1(\dacArea_dac_cnt_3[6] ),
    .A2(net24),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3707_ (.A1(\dacArea_dac_cnt_3[6] ),
    .A2(net24),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3708_ (.A1(_3225_),
    .A2(_3223_),
    .B(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3709_ (.A1(net146),
    .A2(net25),
    .A3(_3227_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3710_ (.A1(_3112_),
    .A2(_3228_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3711_ (.A1(\dacArea_dac_cnt_4[0] ),
    .A2(net26),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3712_ (.A1(\dacArea_dac_cnt_4[0] ),
    .A2(net26),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3713_ (.A1(_3142_),
    .A2(_3229_),
    .A3(_3230_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3714_ (.A1(\dacArea_dac_cnt_4[1] ),
    .A2(net27),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3715_ (.A1(_3230_),
    .A2(_3231_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3716_ (.A1(_3230_),
    .A2(_3231_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3717_ (.A1(_3173_),
    .A2(_3232_),
    .A3(_3233_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3718_ (.I(_3110_),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3719_ (.A1(\dacArea_dac_cnt_4[1] ),
    .A2(net27),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3720_ (.A1(_3235_),
    .A2(_3233_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3721_ (.A1(\dacArea_dac_cnt_4[2] ),
    .A2(net28),
    .A3(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3722_ (.A1(_3234_),
    .A2(_3237_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3723_ (.A1(\dacArea_dac_cnt_4[2] ),
    .A2(net28),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3724_ (.A1(_3236_),
    .A2(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3725_ (.A1(\dacArea_dac_cnt_4[2] ),
    .A2(net28),
    .B(_3239_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3726_ (.A1(\dacArea_dac_cnt_4[3] ),
    .A2(net29),
    .A3(_3240_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3727_ (.A1(_3234_),
    .A2(_3241_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3728_ (.A1(\dacArea_dac_cnt_4[3] ),
    .A2(net29),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3729_ (.A1(\dacArea_dac_cnt_4[3] ),
    .A2(net29),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3730_ (.A1(_3242_),
    .A2(_3240_),
    .B(_3243_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3731_ (.A1(\dacArea_dac_cnt_4[4] ),
    .A2(net30),
    .A3(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3732_ (.A1(_3234_),
    .A2(_3245_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3733_ (.A1(\dacArea_dac_cnt_4[4] ),
    .A2(net30),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3734_ (.A1(\dacArea_dac_cnt_4[4] ),
    .A2(net30),
    .B(_3244_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3735_ (.A1(_3246_),
    .A2(_3247_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3736_ (.A1(\dacArea_dac_cnt_4[5] ),
    .A2(net31),
    .A3(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3737_ (.A1(_3234_),
    .A2(_3249_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3738_ (.A1(\dacArea_dac_cnt_4[5] ),
    .A2(net31),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3739_ (.A1(\dacArea_dac_cnt_4[5] ),
    .A2(net31),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3740_ (.A1(_3250_),
    .A2(_3248_),
    .B(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3741_ (.I(_3252_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3742_ (.A1(\dacArea_dac_cnt_4[6] ),
    .A2(net32),
    .A3(_3253_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3743_ (.A1(_3234_),
    .A2(_3254_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3744_ (.A1(\dacArea_dac_cnt_4[6] ),
    .A2(net32),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3745_ (.A1(\dacArea_dac_cnt_4[6] ),
    .A2(net32),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3746_ (.A1(_3255_),
    .A2(_3253_),
    .B(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3747_ (.A1(net147),
    .A2(net33),
    .A3(_3257_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3748_ (.A1(_3112_),
    .A2(_3258_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3749_ (.A1(\dacArea_dac_cnt_5[0] ),
    .A2(net35),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3750_ (.A1(\dacArea_dac_cnt_5[0] ),
    .A2(net35),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3751_ (.A1(_3142_),
    .A2(_3259_),
    .A3(_3260_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3752_ (.A1(\dacArea_dac_cnt_5[1] ),
    .A2(net36),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3753_ (.A1(_3260_),
    .A2(_3261_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3754_ (.A1(_3260_),
    .A2(_3261_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3755_ (.A1(_3173_),
    .A2(_3262_),
    .A3(_3263_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3756_ (.A1(\dacArea_dac_cnt_5[1] ),
    .A2(net36),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3757_ (.A1(_3264_),
    .A2(_3263_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3758_ (.A1(\dacArea_dac_cnt_5[2] ),
    .A2(net37),
    .A3(_3265_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3759_ (.A1(_3234_),
    .A2(_3266_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3760_ (.A1(\dacArea_dac_cnt_5[2] ),
    .A2(net37),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3761_ (.A1(_3265_),
    .A2(_3267_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3762_ (.A1(\dacArea_dac_cnt_5[2] ),
    .A2(net37),
    .B(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3763_ (.A1(\dacArea_dac_cnt_5[3] ),
    .A2(net38),
    .A3(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3764_ (.A1(_3234_),
    .A2(_3270_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3765_ (.A1(\dacArea_dac_cnt_5[3] ),
    .A2(net38),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3766_ (.A1(\dacArea_dac_cnt_5[3] ),
    .A2(net38),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3767_ (.A1(_3271_),
    .A2(_3269_),
    .B(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3768_ (.A1(\dacArea_dac_cnt_5[4] ),
    .A2(net39),
    .A3(_3273_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3769_ (.A1(_3234_),
    .A2(_3274_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3770_ (.A1(\dacArea_dac_cnt_5[4] ),
    .A2(net39),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3771_ (.A1(\dacArea_dac_cnt_5[4] ),
    .A2(net39),
    .B(_3273_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3772_ (.A1(_3275_),
    .A2(_3276_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3773_ (.A1(\dacArea_dac_cnt_5[5] ),
    .A2(net40),
    .A3(_3277_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3774_ (.A1(_3234_),
    .A2(_3278_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3775_ (.A1(\dacArea_dac_cnt_5[5] ),
    .A2(net40),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3776_ (.A1(_3279_),
    .A2(_3277_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3777_ (.A1(\dacArea_dac_cnt_5[5] ),
    .A2(net40),
    .B(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3778_ (.A1(\dacArea_dac_cnt_5[6] ),
    .A2(net41),
    .A3(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3779_ (.A1(_3234_),
    .A2(_3282_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3780_ (.A1(\dacArea_dac_cnt_5[6] ),
    .A2(net41),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3781_ (.A1(\dacArea_dac_cnt_5[6] ),
    .A2(net41),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3782_ (.A1(_3283_),
    .A2(_3281_),
    .B(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3783_ (.A1(net148),
    .A2(net42),
    .A3(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3784_ (.A1(_3112_),
    .A2(_3286_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3785_ (.A1(\dacArea_dac_cnt_6[0] ),
    .A2(net43),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3786_ (.A1(\dacArea_dac_cnt_6[0] ),
    .A2(net43),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3787_ (.A1(_3142_),
    .A2(_3287_),
    .A3(_3288_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3788_ (.A1(\dacArea_dac_cnt_6[1] ),
    .A2(net44),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3789_ (.A1(_3288_),
    .A2(_3289_),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3790_ (.A1(_3288_),
    .A2(_3289_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3791_ (.A1(_3173_),
    .A2(_3290_),
    .A3(_3291_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3792_ (.I(_3110_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3793_ (.A1(\dacArea_dac_cnt_6[1] ),
    .A2(net44),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3794_ (.A1(_3293_),
    .A2(_3291_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3795_ (.A1(\dacArea_dac_cnt_6[2] ),
    .A2(net46),
    .A3(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3796_ (.A1(_3292_),
    .A2(_3295_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3797_ (.A1(\dacArea_dac_cnt_6[2] ),
    .A2(net46),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3798_ (.A1(_3294_),
    .A2(_3296_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3799_ (.A1(\dacArea_dac_cnt_6[2] ),
    .A2(net46),
    .B(_3297_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3800_ (.A1(\dacArea_dac_cnt_6[3] ),
    .A2(net47),
    .A3(_3298_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3801_ (.A1(_3292_),
    .A2(_3299_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3802_ (.A1(\dacArea_dac_cnt_6[3] ),
    .A2(net47),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3803_ (.A1(\dacArea_dac_cnt_6[3] ),
    .A2(net47),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3804_ (.A1(_3300_),
    .A2(_3298_),
    .B(_3301_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3805_ (.A1(\dacArea_dac_cnt_6[4] ),
    .A2(net48),
    .A3(_3302_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3806_ (.A1(_3292_),
    .A2(_3303_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3807_ (.A1(\dacArea_dac_cnt_6[4] ),
    .A2(net48),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3808_ (.A1(\dacArea_dac_cnt_6[4] ),
    .A2(net48),
    .B(_3302_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3809_ (.A1(_3304_),
    .A2(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3810_ (.A1(\dacArea_dac_cnt_6[5] ),
    .A2(net49),
    .A3(_3306_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3811_ (.A1(_3292_),
    .A2(_3307_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3812_ (.A1(\dacArea_dac_cnt_6[5] ),
    .A2(net49),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3813_ (.A1(_3308_),
    .A2(_3306_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3814_ (.A1(\dacArea_dac_cnt_6[5] ),
    .A2(net49),
    .B(_3309_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3815_ (.A1(\dacArea_dac_cnt_6[6] ),
    .A2(net50),
    .A3(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3816_ (.A1(_3292_),
    .A2(_3311_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3817_ (.A1(\dacArea_dac_cnt_6[6] ),
    .A2(net50),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3818_ (.A1(\dacArea_dac_cnt_6[6] ),
    .A2(net50),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3819_ (.A1(_3312_),
    .A2(_3310_),
    .B(_3313_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3820_ (.A1(net150),
    .A2(net51),
    .A3(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3821_ (.A1(_3112_),
    .A2(_3315_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3822_ (.A1(\dacArea_dac_cnt_7[0] ),
    .A2(net52),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3823_ (.A1(\dacArea_dac_cnt_7[0] ),
    .A2(net52),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3824_ (.A1(_3142_),
    .A2(_3316_),
    .A3(_3317_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3825_ (.A1(\dacArea_dac_cnt_7[1] ),
    .A2(net53),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3826_ (.A1(_3317_),
    .A2(_3318_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3827_ (.A1(_3317_),
    .A2(_3318_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3828_ (.A1(_3173_),
    .A2(_3319_),
    .A3(_3320_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3829_ (.A1(\dacArea_dac_cnt_7[1] ),
    .A2(net53),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3830_ (.A1(_3321_),
    .A2(_3320_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3831_ (.A1(\dacArea_dac_cnt_7[2] ),
    .A2(net54),
    .A3(_3322_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3832_ (.A1(_3292_),
    .A2(_3323_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3833_ (.A1(\dacArea_dac_cnt_7[2] ),
    .A2(net54),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3834_ (.A1(_3322_),
    .A2(_3324_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3835_ (.A1(\dacArea_dac_cnt_7[2] ),
    .A2(net54),
    .B(_3325_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3836_ (.A1(\dacArea_dac_cnt_7[3] ),
    .A2(net55),
    .A3(_3326_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3837_ (.A1(_3292_),
    .A2(_3327_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3838_ (.A1(\dacArea_dac_cnt_7[3] ),
    .A2(net55),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3839_ (.A1(\dacArea_dac_cnt_7[3] ),
    .A2(net55),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3840_ (.A1(_3328_),
    .A2(_3326_),
    .B(_3329_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3841_ (.A1(\dacArea_dac_cnt_7[4] ),
    .A2(net57),
    .A3(_3330_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3842_ (.A1(_3292_),
    .A2(_3331_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3843_ (.A1(\dacArea_dac_cnt_7[4] ),
    .A2(net57),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3844_ (.A1(\dacArea_dac_cnt_7[4] ),
    .A2(net57),
    .B(_3330_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3845_ (.A1(_3332_),
    .A2(_3333_),
    .Z(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3846_ (.A1(\dacArea_dac_cnt_7[5] ),
    .A2(net58),
    .A3(_3334_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3847_ (.A1(_3292_),
    .A2(_3335_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3848_ (.A1(\dacArea_dac_cnt_7[5] ),
    .A2(net58),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3849_ (.A1(_3336_),
    .A2(_3334_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3850_ (.A1(\dacArea_dac_cnt_7[5] ),
    .A2(net58),
    .B(_3337_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3851_ (.A1(\dacArea_dac_cnt_7[6] ),
    .A2(net59),
    .A3(_3338_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3852_ (.A1(_3292_),
    .A2(_3339_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3853_ (.A1(\dacArea_dac_cnt_7[6] ),
    .A2(net59),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3854_ (.A1(\dacArea_dac_cnt_7[6] ),
    .A2(net59),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3855_ (.A1(_3340_),
    .A2(_3338_),
    .B(_3341_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3856_ (.A1(net151),
    .A2(net60),
    .A3(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3857_ (.A1(_3112_),
    .A2(_3343_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3858_ (.I(net99),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3859_ (.A1(net98),
    .A2(net125),
    .A3(net159),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3860_ (.A1(_2989_),
    .A2(_2996_),
    .A3(_3345_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3861_ (.I(_3346_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3862_ (.I(_3346_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3863_ (.A1(_3002_),
    .A2(_3348_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3864_ (.I(_3109_),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3865_ (.A1(_3344_),
    .A2(_3347_),
    .B(_3349_),
    .C(_3350_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3866_ (.I(net110),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3867_ (.A1(_3009_),
    .A2(_3348_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3868_ (.A1(_3351_),
    .A2(_3347_),
    .B(_3352_),
    .C(_3350_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3869_ (.I(net116),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3870_ (.A1(_3013_),
    .A2(_3348_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3871_ (.A1(_3353_),
    .A2(_3347_),
    .B(_3354_),
    .C(_3350_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3872_ (.I(net117),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3873_ (.A1(_3017_),
    .A2(_3348_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3874_ (.A1(_3355_),
    .A2(_3347_),
    .B(_3356_),
    .C(_3350_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3875_ (.I(net118),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3876_ (.A1(_3021_),
    .A2(_3348_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3877_ (.A1(_3357_),
    .A2(_3347_),
    .B(_3358_),
    .C(_3350_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3878_ (.I(net119),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3879_ (.I(_3346_),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3880_ (.A1(_3026_),
    .A2(_3360_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3881_ (.A1(_3359_),
    .A2(_3347_),
    .B(_3361_),
    .C(_3350_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3882_ (.I(net120),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3883_ (.A1(_3030_),
    .A2(_3360_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3884_ (.A1(_3362_),
    .A2(_3347_),
    .B(_3363_),
    .C(_3350_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3885_ (.I(net121),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3886_ (.A1(_3034_),
    .A2(_3360_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3887_ (.A1(_3364_),
    .A2(_3347_),
    .B(_3365_),
    .C(_3350_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3888_ (.I(net122),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3889_ (.A1(_3038_),
    .A2(_3360_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3890_ (.A1(_3366_),
    .A2(_3347_),
    .B(_3367_),
    .C(_3350_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3891_ (.I(net123),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3892_ (.A1(_3042_),
    .A2(_3360_),
    .ZN(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3893_ (.A1(_3368_),
    .A2(_3347_),
    .B(_3369_),
    .C(_3350_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3894_ (.I(net100),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3895_ (.I(_3346_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3896_ (.A1(_3046_),
    .A2(_3360_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3897_ (.I(_3109_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3898_ (.A1(_3370_),
    .A2(_3371_),
    .B(_3372_),
    .C(_3373_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3899_ (.I(net101),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3900_ (.A1(_3050_),
    .A2(_3360_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3901_ (.A1(_3374_),
    .A2(_3371_),
    .B(_3375_),
    .C(_3373_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3902_ (.I(net102),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3903_ (.A1(_3054_),
    .A2(_3360_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3904_ (.A1(_3376_),
    .A2(_3371_),
    .B(_3377_),
    .C(_3373_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3905_ (.I(net103),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3906_ (.A1(_3058_),
    .A2(_3360_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3907_ (.A1(_3378_),
    .A2(_3371_),
    .B(_3379_),
    .C(_3373_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3908_ (.I(net104),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3909_ (.A1(_3062_),
    .A2(_3360_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3910_ (.A1(_3380_),
    .A2(_3371_),
    .B(_3381_),
    .C(_3373_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3911_ (.I(net105),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3912_ (.I(_3346_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3913_ (.A1(_3066_),
    .A2(_3383_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3914_ (.A1(_3382_),
    .A2(_3371_),
    .B(_3384_),
    .C(_3373_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3915_ (.I(net106),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3916_ (.A1(_3070_),
    .A2(_3383_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3917_ (.A1(_3385_),
    .A2(_3371_),
    .B(_3386_),
    .C(_3373_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3918_ (.I(net107),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3919_ (.A1(_3076_),
    .A2(_3383_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3920_ (.A1(_3387_),
    .A2(_3371_),
    .B(_3388_),
    .C(_3373_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3921_ (.I(net108),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3922_ (.A1(_3081_),
    .A2(_3383_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3923_ (.A1(_3389_),
    .A2(_3371_),
    .B(_3390_),
    .C(_3373_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3924_ (.I(net109),
    .ZN(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3925_ (.A1(_3086_),
    .A2(_3383_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3926_ (.A1(_3391_),
    .A2(_3371_),
    .B(_0154_),
    .C(_3373_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3927_ (.I(net111),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3928_ (.A1(_3090_),
    .A2(_3383_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3929_ (.I(_3109_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3930_ (.A1(_0155_),
    .A2(_3348_),
    .B(_0156_),
    .C(_0157_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3931_ (.I(net112),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3932_ (.A1(_3094_),
    .A2(_3383_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3933_ (.A1(_0158_),
    .A2(_3348_),
    .B(_0159_),
    .C(_0157_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3934_ (.I(net113),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3935_ (.A1(_3098_),
    .A2(_3383_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3936_ (.A1(_0160_),
    .A2(_3348_),
    .B(_0161_),
    .C(_0157_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3937_ (.I(net114),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3938_ (.A1(_3102_),
    .A2(_3383_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3939_ (.A1(_0162_),
    .A2(_3348_),
    .B(_0163_),
    .C(_0157_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3940_ (.I(net115),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3941_ (.A1(_3106_),
    .A2(_3383_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3942_ (.A1(_0164_),
    .A2(_3348_),
    .B(_0165_),
    .C(_0157_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3943_ (.I(_3110_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3944_ (.I(\dspArea_regB[0] ),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3945_ (.I(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _3946_ (.A1(_2994_),
    .A2(_2986_),
    .A3(_2990_),
    .A4(_3345_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3947_ (.I(_0169_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3948_ (.I0(_0168_),
    .I1(net99),
    .S(_0170_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3949_ (.A1(_0166_),
    .A2(_0171_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3950_ (.I(\dspArea_regB[1] ),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3951_ (.I(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3952_ (.I(_0173_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3953_ (.I0(_0174_),
    .I1(net110),
    .S(_0170_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3954_ (.A1(_0166_),
    .A2(_0175_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3955_ (.I(\dspArea_regB[2] ),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3956_ (.I(_0176_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3957_ (.I(_0177_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3958_ (.I0(_0178_),
    .I1(net116),
    .S(_0170_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3959_ (.A1(_0166_),
    .A2(_0179_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3960_ (.I(\dspArea_regB[3] ),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3961_ (.I(_0180_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3962_ (.I(_0181_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3963_ (.I(_0182_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3964_ (.I(_0183_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3965_ (.I0(_0184_),
    .I1(net117),
    .S(_0170_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3966_ (.A1(_0166_),
    .A2(_0185_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3967_ (.I(\dspArea_regB[4] ),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3968_ (.I(_0186_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3969_ (.I(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3970_ (.I(_0188_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3971_ (.I(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3972_ (.I0(_0190_),
    .I1(net118),
    .S(_0170_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3973_ (.A1(_0166_),
    .A2(_0191_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3974_ (.I(\dspArea_regB[5] ),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3975_ (.I(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3976_ (.I0(_0193_),
    .I1(net119),
    .S(_0170_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3977_ (.A1(_0166_),
    .A2(_0194_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3978_ (.I(\dspArea_regB[6] ),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3979_ (.I(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3980_ (.I(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3981_ (.I(_0197_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3982_ (.I0(_0198_),
    .I1(net120),
    .S(_0170_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3983_ (.A1(_0166_),
    .A2(_0199_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3984_ (.I(\dspArea_regB[7] ),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3985_ (.I(_0200_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3986_ (.I(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3987_ (.I(_0202_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3988_ (.I0(_0203_),
    .I1(net121),
    .S(_0170_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3989_ (.A1(_0166_),
    .A2(_0204_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3990_ (.I(\dspArea_regB[8] ),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3991_ (.I(_0205_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3992_ (.I(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3993_ (.I0(_0207_),
    .I1(net122),
    .S(_0170_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3994_ (.A1(_0166_),
    .A2(_0208_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3995_ (.I(\dspArea_regB[9] ),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3996_ (.I(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3997_ (.I(_0210_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3998_ (.I(_0211_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3999_ (.I(_0212_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4000_ (.I0(_0213_),
    .I1(net123),
    .S(_0170_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4001_ (.A1(_0166_),
    .A2(_0214_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4002_ (.I(_3110_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4003_ (.I(\dspArea_regB[10] ),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4004_ (.I(_0216_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4005_ (.I(_0217_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4006_ (.I(_0218_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4007_ (.I0(_0219_),
    .I1(net100),
    .S(_0169_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4008_ (.A1(_0215_),
    .A2(_0220_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4009_ (.I(\dspArea_regB[11] ),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4010_ (.I(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4011_ (.I(_0222_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4012_ (.I0(_0223_),
    .I1(net101),
    .S(_0169_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4013_ (.A1(_0215_),
    .A2(_0224_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4014_ (.I(\dspArea_regB[12] ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4015_ (.I(_0225_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4016_ (.I(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4017_ (.I(_0227_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4018_ (.I(_0228_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4019_ (.I0(_0229_),
    .I1(net102),
    .S(_0169_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4020_ (.A1(_0215_),
    .A2(_0230_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4021_ (.I(\dspArea_regB[13] ),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4022_ (.I(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4023_ (.I(_0232_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4024_ (.I(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4025_ (.I0(_0234_),
    .I1(net103),
    .S(_0169_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4026_ (.A1(_0215_),
    .A2(_0235_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4027_ (.I(\dspArea_regB[14] ),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4028_ (.I(_0236_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4029_ (.I(_0237_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4030_ (.I0(_0238_),
    .I1(net104),
    .S(_0169_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4031_ (.A1(_0215_),
    .A2(_0239_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4032_ (.I(\dspArea_regB[15] ),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4033_ (.I(_0240_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4034_ (.I(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4035_ (.I(_0242_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4036_ (.I(_0243_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4037_ (.I0(_0244_),
    .I1(net105),
    .S(_0169_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4038_ (.A1(_0215_),
    .A2(_0245_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4039_ (.A1(_2985_),
    .A2(_2995_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4040_ (.I(_0246_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4041_ (.A1(net98),
    .A2(net159),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4042_ (.A1(net125),
    .A2(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4043_ (.A1(_2982_),
    .A2(_2997_),
    .A3(_0247_),
    .A4(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4044_ (.A1(_0168_),
    .A2(_3002_),
    .A3(_0250_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4045_ (.A1(\dspArea_regP[0] ),
    .A2(_0251_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4046_ (.A1(_0215_),
    .A2(_0252_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4047_ (.A1(\dspArea_regP[0] ),
    .A2(_0168_),
    .A3(_3002_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4048_ (.A1(_0168_),
    .A2(_3009_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4049_ (.A1(\dspArea_regP[1] ),
    .A2(_0254_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4050_ (.A1(_0174_),
    .A2(_3002_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4051_ (.A1(_0255_),
    .A2(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4052_ (.A1(_0253_),
    .A2(_0257_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4053_ (.I(_0250_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4054_ (.I0(\dspArea_regP[1] ),
    .I1(_0258_),
    .S(_0259_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4055_ (.A1(_0215_),
    .A2(_0260_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4056_ (.A1(_0253_),
    .A2(_0257_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4057_ (.A1(_0168_),
    .A2(_3013_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4058_ (.A1(\dspArea_regP[2] ),
    .A2(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4059_ (.A1(_0174_),
    .A2(_3009_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4060_ (.A1(_0263_),
    .A2(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4061_ (.A1(\dspArea_regP[1] ),
    .A2(_0254_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4062_ (.A1(_0255_),
    .A2(_0256_),
    .B(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4063_ (.A1(_0265_),
    .A2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4064_ (.A1(_0178_),
    .A2(_3002_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4065_ (.A1(_0268_),
    .A2(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4066_ (.A1(_0261_),
    .A2(_0270_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4067_ (.I0(\dspArea_regP[2] ),
    .I1(_0271_),
    .S(_0259_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4068_ (.A1(_0215_),
    .A2(_0272_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4069_ (.A1(_0261_),
    .A2(_0270_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4070_ (.A1(_0174_),
    .A2(_3013_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4071_ (.A1(_0168_),
    .A2(_3017_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4072_ (.A1(\dspArea_regP[3] ),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4073_ (.A1(_0274_),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4074_ (.A1(\dspArea_regP[2] ),
    .A2(_0262_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4075_ (.A1(_0263_),
    .A2(_0264_),
    .B(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4076_ (.A1(_0277_),
    .A2(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4077_ (.A1(_0178_),
    .A2(_3009_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4078_ (.A1(_0184_),
    .A2(_3002_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4079_ (.A1(_0184_),
    .A2(_3008_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4080_ (.A1(_0269_),
    .A2(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4081_ (.A1(_0281_),
    .A2(_0282_),
    .B(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4082_ (.A1(_0280_),
    .A2(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4083_ (.I(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4084_ (.I(_0265_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4085_ (.A1(_0288_),
    .A2(_0267_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4086_ (.A1(_0178_),
    .A2(_3002_),
    .A3(_0268_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4087_ (.A1(_0289_),
    .A2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4088_ (.A1(_0287_),
    .A2(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4089_ (.A1(_0273_),
    .A2(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4090_ (.I0(\dspArea_regP[3] ),
    .I1(_0293_),
    .S(_0259_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4091_ (.A1(_0215_),
    .A2(_0294_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4092_ (.I(\dspArea_regP[4] ),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4093_ (.A1(_2998_),
    .A2(_0249_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4094_ (.I(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4095_ (.A1(_2998_),
    .A2(_0249_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4096_ (.I(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4097_ (.A1(_0178_),
    .A2(_3012_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4098_ (.A1(_0283_),
    .A2(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4099_ (.A1(_0190_),
    .A2(_3001_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4100_ (.A1(_0301_),
    .A2(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4101_ (.I(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4102_ (.A1(_0174_),
    .A2(_3017_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4103_ (.A1(_0168_),
    .A2(_3020_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4104_ (.A1(\dspArea_regP[4] ),
    .A2(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4105_ (.A1(_0305_),
    .A2(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4106_ (.A1(\dspArea_regP[3] ),
    .A2(_0275_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4107_ (.A1(_0274_),
    .A2(_0276_),
    .B(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4108_ (.A1(_0304_),
    .A2(_0308_),
    .A3(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4109_ (.A1(_0277_),
    .A2(_0279_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4110_ (.I(_0285_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4111_ (.A1(_0280_),
    .A2(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4112_ (.A1(_0312_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4113_ (.A1(_0284_),
    .A2(_0311_),
    .A3(_0315_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4114_ (.A1(_0287_),
    .A2(_0291_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4115_ (.A1(_0273_),
    .A2(_0292_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4116_ (.A1(_0317_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4117_ (.A1(_0316_),
    .A2(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4118_ (.A1(_0316_),
    .A2(_0319_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4119_ (.A1(_0299_),
    .A2(_0320_),
    .A3(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4120_ (.A1(_0295_),
    .A2(_0297_),
    .B(_0322_),
    .C(_0157_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4121_ (.A1(_0318_),
    .A2(_0316_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4122_ (.A1(_0317_),
    .A2(_0316_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4123_ (.A1(_0184_),
    .A2(_3013_),
    .A3(_0281_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4124_ (.A1(_0190_),
    .A2(_3001_),
    .A3(_0301_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4125_ (.A1(_0325_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4126_ (.A1(_0193_),
    .A2(_3000_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4127_ (.A1(_0327_),
    .A2(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4128_ (.I(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4129_ (.A1(_0190_),
    .A2(_3008_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4130_ (.A1(_0182_),
    .A2(_3012_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4131_ (.A1(_0177_),
    .A2(_3016_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4132_ (.A1(_0332_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4133_ (.A1(_0331_),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4134_ (.I(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4135_ (.A1(_0174_),
    .A2(_3020_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4136_ (.A1(_0167_),
    .A2(_3025_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4137_ (.A1(\dspArea_regP[5] ),
    .A2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4138_ (.A1(_0337_),
    .A2(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4139_ (.A1(\dspArea_regP[4] ),
    .A2(_0306_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4140_ (.A1(_0305_),
    .A2(_0307_),
    .B(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4141_ (.A1(_0336_),
    .A2(_0340_),
    .A3(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4142_ (.A1(_0308_),
    .A2(_0310_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4143_ (.A1(_0308_),
    .A2(_0310_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4144_ (.A1(_0304_),
    .A2(_0344_),
    .B(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4145_ (.A1(_0330_),
    .A2(_0343_),
    .A3(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4146_ (.A1(_0312_),
    .A2(_0314_),
    .A3(_0311_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4147_ (.A1(_0312_),
    .A2(_0314_),
    .B(_0311_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4148_ (.A1(_0284_),
    .A2(_0348_),
    .B(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4149_ (.A1(_0347_),
    .A2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4150_ (.A1(_0324_),
    .A2(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4151_ (.A1(_0323_),
    .A2(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4152_ (.A1(\dspArea_regP[5] ),
    .A2(_0299_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4153_ (.A1(_0299_),
    .A2(_0353_),
    .B(_0354_),
    .C(_0157_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4154_ (.I(_3110_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4155_ (.A1(_0323_),
    .A2(_0352_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4156_ (.A1(_0325_),
    .A2(_0326_),
    .B(_0328_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4157_ (.A1(_0184_),
    .A2(_3017_),
    .A3(_0300_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4158_ (.A1(_0190_),
    .A2(_3008_),
    .A3(_0334_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4159_ (.A1(_0358_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4160_ (.A1(_0193_),
    .A2(_3008_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4161_ (.A1(_0198_),
    .A2(_3000_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4162_ (.A1(_0361_),
    .A2(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4163_ (.I(_0195_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4164_ (.A1(_0364_),
    .A2(_3007_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4165_ (.A1(_0328_),
    .A2(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4166_ (.A1(_0363_),
    .A2(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4167_ (.A1(_0360_),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4168_ (.I(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4169_ (.A1(_0187_),
    .A2(_3012_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4170_ (.A1(_0181_),
    .A2(_3015_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4171_ (.A1(_0176_),
    .A2(_3019_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4172_ (.A1(_0371_),
    .A2(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4173_ (.A1(_0370_),
    .A2(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4174_ (.I(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4175_ (.A1(\dspArea_regP[5] ),
    .A2(_0168_),
    .A3(_3025_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4176_ (.I(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4177_ (.A1(_0337_),
    .A2(_0339_),
    .B(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4178_ (.A1(_0174_),
    .A2(_3026_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4179_ (.A1(_0168_),
    .A2(_3029_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4180_ (.A1(\dspArea_regP[6] ),
    .A2(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4181_ (.A1(_0379_),
    .A2(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4182_ (.A1(_0375_),
    .A2(_0378_),
    .A3(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4183_ (.A1(_0340_),
    .A2(_0342_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4184_ (.A1(_0340_),
    .A2(_0342_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4185_ (.A1(_0336_),
    .A2(_0384_),
    .B(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4186_ (.A1(_0383_),
    .A2(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4187_ (.A1(_0369_),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4188_ (.A1(_0343_),
    .A2(_0346_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4189_ (.A1(_0343_),
    .A2(_0346_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4190_ (.A1(_0330_),
    .A2(_0389_),
    .B(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4191_ (.A1(_0357_),
    .A2(_0388_),
    .A3(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4192_ (.A1(_0347_),
    .A2(_0350_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4193_ (.A1(_0324_),
    .A2(_0351_),
    .B(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4194_ (.A1(_0392_),
    .A2(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4195_ (.A1(_0356_),
    .A2(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4196_ (.I0(\dspArea_regP[6] ),
    .I1(_0396_),
    .S(_0259_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4197_ (.A1(_0355_),
    .A2(_0397_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4198_ (.A1(_0356_),
    .A2(_0395_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4199_ (.A1(_0347_),
    .A2(_0350_),
    .A3(_0392_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4200_ (.A1(_0360_),
    .A2(_0367_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4201_ (.A1(_0183_),
    .A2(_3021_),
    .A3(_0333_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4202_ (.A1(_0189_),
    .A2(_3012_),
    .A3(_0373_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4203_ (.A1(_0401_),
    .A2(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4204_ (.I(_0200_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4205_ (.A1(_0404_),
    .A2(_3000_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4206_ (.I(_0192_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4207_ (.A1(_0406_),
    .A2(_3011_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4208_ (.A1(_0365_),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4209_ (.A1(_0405_),
    .A2(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4210_ (.A1(_0403_),
    .A2(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4211_ (.A1(_0366_),
    .A2(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4212_ (.A1(_0188_),
    .A2(_3016_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4213_ (.A1(_0181_),
    .A2(_3019_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4214_ (.A1(_0177_),
    .A2(_3024_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4215_ (.A1(_0413_),
    .A2(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4216_ (.A1(_0412_),
    .A2(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4217_ (.I(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4218_ (.A1(_0174_),
    .A2(_3030_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4219_ (.A1(_0167_),
    .A2(_3033_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4220_ (.A1(\dspArea_regP[7] ),
    .A2(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4221_ (.A1(_0418_),
    .A2(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4222_ (.A1(\dspArea_regP[6] ),
    .A2(_0380_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4223_ (.A1(_0379_),
    .A2(_0381_),
    .B(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4224_ (.A1(_0417_),
    .A2(_0421_),
    .A3(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4225_ (.A1(_0378_),
    .A2(_0382_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4226_ (.A1(_0378_),
    .A2(_0382_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4227_ (.A1(_0375_),
    .A2(_0425_),
    .B(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4228_ (.A1(_0411_),
    .A2(_0424_),
    .A3(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4229_ (.A1(_0383_),
    .A2(_0386_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4230_ (.A1(_0383_),
    .A2(_0386_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4231_ (.A1(_0369_),
    .A2(_0429_),
    .B(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4232_ (.A1(_0428_),
    .A2(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4233_ (.A1(_0400_),
    .A2(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4234_ (.A1(_0388_),
    .A2(_0391_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4235_ (.A1(_0388_),
    .A2(_0391_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4236_ (.A1(_0357_),
    .A2(_0434_),
    .B(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4237_ (.A1(_0399_),
    .A2(_0433_),
    .A3(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4238_ (.A1(_0324_),
    .A2(_0351_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4239_ (.A1(_0438_),
    .A2(_0392_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4240_ (.A1(_0398_),
    .A2(_0437_),
    .A3(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4241_ (.I(_0250_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4242_ (.I0(\dspArea_regP[7] ),
    .I1(_0440_),
    .S(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4243_ (.A1(_0355_),
    .A2(_0442_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4244_ (.A1(_0437_),
    .A2(_0439_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4245_ (.A1(_0437_),
    .A2(_0439_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4246_ (.A1(_0398_),
    .A2(_0443_),
    .B(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4247_ (.I(_0403_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4248_ (.A1(_0446_),
    .A2(_0409_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4249_ (.A1(_0366_),
    .A2(_0410_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4250_ (.A1(_0447_),
    .A2(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4251_ (.A1(_0207_),
    .A2(_3001_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4252_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4253_ (.A1(_0364_),
    .A2(_3011_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4254_ (.A1(_0361_),
    .A2(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4255_ (.A1(_0203_),
    .A2(_3000_),
    .A3(_0408_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4256_ (.A1(_0453_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4257_ (.A1(_0183_),
    .A2(_3025_),
    .A3(_0372_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4258_ (.A1(_0189_),
    .A2(_3016_),
    .A3(_0415_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4259_ (.A1(_0456_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4260_ (.A1(_0201_),
    .A2(_3008_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4261_ (.A1(_0406_),
    .A2(_3015_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4262_ (.A1(_0452_),
    .A2(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4263_ (.A1(_0459_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4264_ (.A1(_0458_),
    .A2(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4265_ (.A1(_0455_),
    .A2(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4266_ (.A1(_0187_),
    .A2(_3020_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4267_ (.A1(_0181_),
    .A2(_3024_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4268_ (.A1(_0176_),
    .A2(_3028_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4269_ (.A1(_0466_),
    .A2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4270_ (.A1(_0465_),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4271_ (.I(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4272_ (.A1(_0173_),
    .A2(_3033_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4273_ (.A1(_0167_),
    .A2(_3036_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4274_ (.A1(\dspArea_regP[8] ),
    .A2(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4275_ (.A1(_0471_),
    .A2(_0473_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4276_ (.A1(\dspArea_regP[7] ),
    .A2(_0419_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4277_ (.A1(_0418_),
    .A2(_0420_),
    .B(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4278_ (.A1(_0470_),
    .A2(_0474_),
    .A3(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4279_ (.A1(_0421_),
    .A2(_0423_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4280_ (.A1(_0421_),
    .A2(_0423_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4281_ (.A1(_0417_),
    .A2(_0478_),
    .B(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4282_ (.A1(_0477_),
    .A2(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4283_ (.A1(_0464_),
    .A2(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4284_ (.A1(_0424_),
    .A2(_0427_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4285_ (.A1(_0424_),
    .A2(_0427_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4286_ (.A1(_0411_),
    .A2(_0483_),
    .B(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4287_ (.A1(_0482_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4288_ (.A1(_0451_),
    .A2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4289_ (.A1(_0368_),
    .A2(_0387_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4290_ (.A1(_0430_),
    .A2(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4291_ (.A1(_0360_),
    .A2(_0367_),
    .A3(_0432_),
    .B1(_0489_),
    .B2(_0428_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4292_ (.A1(_0487_),
    .A2(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4293_ (.A1(_0433_),
    .A2(_0436_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4294_ (.A1(_0433_),
    .A2(_0436_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4295_ (.A1(_0399_),
    .A2(_0492_),
    .B(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4296_ (.A1(_0491_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4297_ (.A1(_0445_),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4298_ (.A1(\dspArea_regP[8] ),
    .A2(_0299_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4299_ (.A1(_0299_),
    .A2(_0496_),
    .B(_0497_),
    .C(_0157_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4300_ (.A1(_0445_),
    .A2(_0495_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4301_ (.A1(_0399_),
    .A2(_0492_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4302_ (.A1(_0499_),
    .A2(_0491_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4303_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4304_ (.I(_0458_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4305_ (.A1(_0502_),
    .A2(_0462_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4306_ (.A1(_0455_),
    .A2(_0463_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4307_ (.A1(_0503_),
    .A2(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4308_ (.A1(_0207_),
    .A2(_3008_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4309_ (.A1(_0213_),
    .A2(_3001_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4310_ (.A1(_0505_),
    .A2(_0506_),
    .A3(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4311_ (.A1(_0196_),
    .A2(_3015_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4312_ (.A1(_0407_),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4313_ (.A1(_0203_),
    .A2(_3009_),
    .A3(_0461_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4314_ (.A1(_0510_),
    .A2(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4315_ (.A1(_0184_),
    .A2(_3030_),
    .A3(_0414_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4316_ (.A1(_0189_),
    .A2(_3021_),
    .A3(_0468_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4317_ (.A1(_0513_),
    .A2(_0514_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4318_ (.A1(_0201_),
    .A2(_3012_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4319_ (.A1(_0193_),
    .A2(_3020_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4320_ (.A1(_0509_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4321_ (.A1(_0516_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4322_ (.A1(_0515_),
    .A2(_0519_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4323_ (.A1(_0512_),
    .A2(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4324_ (.A1(_0188_),
    .A2(_3025_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4325_ (.A1(_0181_),
    .A2(_3029_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4326_ (.A1(_0177_),
    .A2(_3032_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4327_ (.A1(_0523_),
    .A2(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4328_ (.A1(_0522_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4329_ (.I(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4330_ (.A1(_0172_),
    .A2(_3037_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4331_ (.I(\dspArea_regB[0] ),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4332_ (.A1(_0529_),
    .A2(_3040_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4333_ (.A1(\dspArea_regP[9] ),
    .A2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4334_ (.A1(_0528_),
    .A2(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4335_ (.A1(\dspArea_regP[8] ),
    .A2(_0472_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4336_ (.A1(_0471_),
    .A2(_0473_),
    .B(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4337_ (.A1(_0532_),
    .A2(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4338_ (.A1(_0527_),
    .A2(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4339_ (.A1(_0474_),
    .A2(_0476_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4340_ (.A1(_0474_),
    .A2(_0476_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4341_ (.A1(_0470_),
    .A2(_0537_),
    .B(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4342_ (.A1(_0536_),
    .A2(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4343_ (.A1(_0521_),
    .A2(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4344_ (.A1(_0477_),
    .A2(_0480_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4345_ (.A1(_0464_),
    .A2(_0481_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4346_ (.A1(_0542_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4347_ (.A1(_0508_),
    .A2(_0541_),
    .A3(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4348_ (.A1(_0482_),
    .A2(_0485_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4349_ (.A1(_0451_),
    .A2(_0486_),
    .B(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4350_ (.A1(_0545_),
    .A2(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4351_ (.A1(_0501_),
    .A2(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4352_ (.A1(_0451_),
    .A2(_0486_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4353_ (.A1(_0550_),
    .A2(_0490_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4354_ (.A1(_0493_),
    .A2(_0491_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4355_ (.A1(_0551_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4356_ (.A1(_0549_),
    .A2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4357_ (.A1(_0498_),
    .A2(_0500_),
    .B(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4358_ (.A1(_0498_),
    .A2(_0500_),
    .A3(_0554_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4359_ (.A1(_0555_),
    .A2(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4360_ (.I0(\dspArea_regP[9] ),
    .I1(_0557_),
    .S(_0441_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4361_ (.A1(_0355_),
    .A2(_0558_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4362_ (.A1(_0549_),
    .A2(_0552_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4363_ (.A1(_0555_),
    .A2(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4364_ (.A1(_0551_),
    .A2(_0549_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4365_ (.A1(_0545_),
    .A2(_0547_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4366_ (.A1(_0501_),
    .A2(_0548_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4367_ (.A1(_0562_),
    .A2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4368_ (.A1(_0506_),
    .A2(_0507_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4369_ (.A1(_0211_),
    .A2(_3007_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4370_ (.A1(_0450_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4371_ (.A1(_0505_),
    .A2(_0565_),
    .A3(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4372_ (.I(_0515_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4373_ (.A1(_0569_),
    .A2(_0519_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4374_ (.A1(_0512_),
    .A2(_0520_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4375_ (.A1(_0570_),
    .A2(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4376_ (.A1(_0207_),
    .A2(_3012_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4377_ (.A1(_0566_),
    .A2(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4378_ (.A1(_0219_),
    .A2(_3001_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4379_ (.A1(_0574_),
    .A2(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4380_ (.A1(_0567_),
    .A2(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4381_ (.A1(_0572_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4382_ (.A1(_0198_),
    .A2(_3021_),
    .A3(_0460_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4383_ (.A1(_0203_),
    .A2(_3013_),
    .A3(_0518_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4384_ (.A1(_0579_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4385_ (.A1(_0182_),
    .A2(_3033_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4386_ (.A1(_0467_),
    .A2(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4387_ (.A1(_0190_),
    .A2(_3026_),
    .A3(_0525_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4388_ (.A1(_0583_),
    .A2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4389_ (.A1(_0201_),
    .A2(_3016_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4390_ (.A1(_0196_),
    .A2(_3020_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4391_ (.A1(_0193_),
    .A2(_3025_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4392_ (.A1(_0587_),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4393_ (.A1(_0586_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4394_ (.A1(_0585_),
    .A2(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4395_ (.A1(_0581_),
    .A2(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4396_ (.A1(_0187_),
    .A2(_3029_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4397_ (.A1(_0178_),
    .A2(_3037_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4398_ (.A1(_0582_),
    .A2(_0593_),
    .A3(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4399_ (.A1(_0174_),
    .A2(_3041_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4400_ (.A1(_0167_),
    .A2(_3044_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4401_ (.A1(\dspArea_regP[10] ),
    .A2(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4402_ (.A1(_0596_),
    .A2(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4403_ (.A1(\dspArea_regP[9] ),
    .A2(_0530_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4404_ (.A1(_0528_),
    .A2(_0531_),
    .B(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4405_ (.A1(_0595_),
    .A2(_0599_),
    .A3(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4406_ (.A1(_0532_),
    .A2(_0534_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4407_ (.A1(_0532_),
    .A2(_0534_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4408_ (.A1(_0527_),
    .A2(_0603_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4409_ (.A1(_0602_),
    .A2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4410_ (.A1(_0592_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4411_ (.A1(_0536_),
    .A2(_0539_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4412_ (.A1(_0521_),
    .A2(_0540_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4413_ (.A1(_0608_),
    .A2(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4414_ (.A1(_0578_),
    .A2(_0607_),
    .A3(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4415_ (.A1(_0542_),
    .A2(_0543_),
    .A3(_0541_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4416_ (.A1(_0542_),
    .A2(_0543_),
    .B(_0541_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4417_ (.A1(_0508_),
    .A2(_0612_),
    .B(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4418_ (.A1(_0611_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4419_ (.A1(_0568_),
    .A2(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4420_ (.A1(_0561_),
    .A2(_0564_),
    .A3(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4421_ (.I(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4422_ (.A1(_0560_),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4423_ (.I0(\dspArea_regP[10] ),
    .I1(_0619_),
    .S(_0441_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4424_ (.A1(_0355_),
    .A2(_0620_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4425_ (.A1(\dspArea_regP[11] ),
    .A2(_0259_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4426_ (.A1(_0562_),
    .A2(_0563_),
    .A3(_0616_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4427_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0616_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4428_ (.A1(_0561_),
    .A2(_0622_),
    .A3(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4429_ (.A1(_0560_),
    .A2(_0617_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4430_ (.A1(_0624_),
    .A2(_0625_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4431_ (.A1(_0572_),
    .A2(_0577_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4432_ (.I(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4433_ (.A1(_0567_),
    .A2(_0576_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4434_ (.I(_0585_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4435_ (.A1(_0630_),
    .A2(_0590_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4436_ (.A1(_0581_),
    .A2(_0591_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4437_ (.A1(_0631_),
    .A2(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4438_ (.I(_0217_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4439_ (.A1(_0634_),
    .A2(_3008_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4440_ (.A1(_0210_),
    .A2(_3011_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4441_ (.A1(_0206_),
    .A2(_3015_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4442_ (.A1(_0636_),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4443_ (.A1(_0635_),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4444_ (.A1(_0506_),
    .A2(_0636_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4445_ (.A1(_0219_),
    .A2(_3000_),
    .A3(_0574_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4446_ (.A1(_0640_),
    .A2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4447_ (.A1(_0639_),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4448_ (.A1(_0223_),
    .A2(_3001_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4449_ (.A1(_0643_),
    .A2(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4450_ (.I(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4451_ (.A1(_0629_),
    .A2(_0633_),
    .A3(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4452_ (.A1(_0198_),
    .A2(_3026_),
    .A3(_0517_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4453_ (.A1(_0203_),
    .A2(_3016_),
    .A3(_0589_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4454_ (.A1(_0648_),
    .A2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4455_ (.A1(_0582_),
    .A2(_0594_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4456_ (.A1(_0182_),
    .A2(_0178_),
    .A3(_3037_),
    .A4(_3033_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4457_ (.I(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4458_ (.A1(_0593_),
    .A2(_0651_),
    .B(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4459_ (.A1(_0404_),
    .A2(_3020_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4460_ (.A1(_0364_),
    .A2(_3024_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4461_ (.A1(_0192_),
    .A2(_3028_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4462_ (.A1(_0656_),
    .A2(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4463_ (.A1(_0655_),
    .A2(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4464_ (.A1(_0654_),
    .A2(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4465_ (.A1(_0650_),
    .A2(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4466_ (.A1(_0182_),
    .A2(_3037_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4467_ (.A1(_0187_),
    .A2(_3033_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4468_ (.A1(_0178_),
    .A2(_3041_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4469_ (.A1(_0662_),
    .A2(_0663_),
    .A3(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4470_ (.I(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4471_ (.A1(_0174_),
    .A2(_3045_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4472_ (.A1(_0167_),
    .A2(_3049_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4473_ (.A1(\dspArea_regP[11] ),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4474_ (.A1(_0667_),
    .A2(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4475_ (.A1(\dspArea_regP[10] ),
    .A2(_0597_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4476_ (.A1(_0596_),
    .A2(_0598_),
    .B(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4477_ (.A1(_0666_),
    .A2(_0670_),
    .A3(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4478_ (.I(_0595_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4479_ (.A1(_0599_),
    .A2(_0601_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4480_ (.A1(_0599_),
    .A2(_0601_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4481_ (.A1(_0674_),
    .A2(_0675_),
    .B(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4482_ (.A1(_0673_),
    .A2(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4483_ (.A1(_0661_),
    .A2(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4484_ (.A1(_0526_),
    .A2(_0535_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4485_ (.A1(_0604_),
    .A2(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4486_ (.A1(_0602_),
    .A2(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4487_ (.A1(_0592_),
    .A2(_0606_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4488_ (.A1(_0682_),
    .A2(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4489_ (.A1(_0647_),
    .A2(_0679_),
    .A3(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4490_ (.A1(_0608_),
    .A2(_0609_),
    .A3(_0607_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4491_ (.A1(_0608_),
    .A2(_0609_),
    .B(_0607_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4492_ (.A1(_0578_),
    .A2(_0686_),
    .B(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4493_ (.A1(_0628_),
    .A2(_0685_),
    .A3(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4494_ (.A1(_0611_),
    .A2(_0614_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4495_ (.A1(_0568_),
    .A2(_0615_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4496_ (.A1(_0690_),
    .A2(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4497_ (.A1(_0689_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4498_ (.A1(_0623_),
    .A2(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4499_ (.A1(_0626_),
    .A2(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4500_ (.A1(_0626_),
    .A2(_0694_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4501_ (.A1(_0297_),
    .A2(_0695_),
    .A3(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4502_ (.A1(_3173_),
    .A2(_0621_),
    .A3(_0697_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4503_ (.A1(_0445_),
    .A2(_0495_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4504_ (.A1(_0499_),
    .A2(_0491_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4505_ (.I(_0549_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4506_ (.A1(_0700_),
    .A2(_0553_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4507_ (.A1(_0700_),
    .A2(_0553_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4508_ (.A1(_0698_),
    .A2(_0699_),
    .B(_0701_),
    .C(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4509_ (.I(_0559_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4510_ (.A1(_0623_),
    .A2(_0693_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4511_ (.A1(_0623_),
    .A2(_0693_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4512_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0705_),
    .B2(_0706_),
    .C(_0617_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4513_ (.I(_0693_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4514_ (.A1(_0623_),
    .A2(_0624_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4515_ (.A1(_0708_),
    .A2(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4516_ (.A1(_0707_),
    .A2(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4517_ (.I(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4518_ (.I(_0689_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4519_ (.A1(_0685_),
    .A2(_0688_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4520_ (.A1(_0685_),
    .A2(_0688_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4521_ (.A1(_0628_),
    .A2(_0714_),
    .B(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4522_ (.A1(_0633_),
    .A2(_0646_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4523_ (.A1(_0633_),
    .A2(_0646_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4524_ (.A1(_0629_),
    .A2(_0718_),
    .A3(_0717_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4525_ (.A1(_0717_),
    .A2(_0719_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4526_ (.I(_0642_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4527_ (.A1(_0639_),
    .A2(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4528_ (.A1(_0223_),
    .A2(_3001_),
    .A3(_0643_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4529_ (.A1(_0722_),
    .A2(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4530_ (.I(_0659_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4531_ (.A1(_0654_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4532_ (.A1(_0650_),
    .A2(_0660_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4533_ (.A1(_0726_),
    .A2(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4534_ (.A1(_0223_),
    .A2(_3008_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4535_ (.A1(_0227_),
    .A2(_3000_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4536_ (.A1(_0729_),
    .A2(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4537_ (.A1(_0217_),
    .A2(_3012_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4538_ (.A1(_0210_),
    .A2(_3015_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4539_ (.A1(_0206_),
    .A2(_3019_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4540_ (.A1(_0733_),
    .A2(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4541_ (.A1(_0732_),
    .A2(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4542_ (.A1(_0212_),
    .A2(_3016_),
    .A3(_0573_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4543_ (.A1(_0218_),
    .A2(_3007_),
    .A3(_0638_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4544_ (.A1(_0737_),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4545_ (.A1(_0736_),
    .A2(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4546_ (.A1(_0731_),
    .A2(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4547_ (.A1(_0728_),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4548_ (.A1(_0724_),
    .A2(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4549_ (.A1(_0198_),
    .A2(_3030_),
    .A3(_0588_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4550_ (.A1(_0655_),
    .A2(_0658_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4551_ (.A1(_0744_),
    .A2(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4552_ (.A1(_0662_),
    .A2(_0664_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4553_ (.A1(_0182_),
    .A2(_0178_),
    .A3(_3041_),
    .A4(_3037_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4554_ (.I(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4555_ (.A1(_0663_),
    .A2(_0747_),
    .B(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4556_ (.A1(_0200_),
    .A2(_3025_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4557_ (.A1(_0364_),
    .A2(_3029_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4558_ (.A1(_0192_),
    .A2(_3032_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4559_ (.A1(_0752_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4560_ (.A1(_0751_),
    .A2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4561_ (.A1(_0750_),
    .A2(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4562_ (.A1(_0746_),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4563_ (.A1(_0181_),
    .A2(_3040_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4564_ (.A1(_0186_),
    .A2(_3036_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4565_ (.A1(_0177_),
    .A2(_3045_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4566_ (.A1(_0758_),
    .A2(_0759_),
    .A3(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4567_ (.I(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4568_ (.A1(_0173_),
    .A2(_3049_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4569_ (.A1(_0167_),
    .A2(_3053_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4570_ (.A1(\dspArea_regP[12] ),
    .A2(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4571_ (.A1(_0763_),
    .A2(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4572_ (.A1(\dspArea_regP[11] ),
    .A2(_0668_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4573_ (.A1(_0667_),
    .A2(_0669_),
    .B(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4574_ (.A1(_0762_),
    .A2(_0766_),
    .A3(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4575_ (.A1(_0670_),
    .A2(_0672_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4576_ (.A1(_0670_),
    .A2(_0672_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4577_ (.A1(_0666_),
    .A2(_0770_),
    .B(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4578_ (.A1(_0769_),
    .A2(_0772_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4579_ (.A1(_0757_),
    .A2(_0773_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4580_ (.A1(_0673_),
    .A2(_0677_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4581_ (.A1(_0661_),
    .A2(_0678_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4582_ (.A1(_0775_),
    .A2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4583_ (.A1(_0743_),
    .A2(_0774_),
    .A3(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4584_ (.A1(_0682_),
    .A2(_0683_),
    .A3(_0679_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4585_ (.A1(_0682_),
    .A2(_0683_),
    .B(_0679_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4586_ (.A1(_0647_),
    .A2(_0779_),
    .B(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4587_ (.A1(_0778_),
    .A2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4588_ (.A1(_0716_),
    .A2(_0720_),
    .A3(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4589_ (.A1(_0713_),
    .A2(_0692_),
    .B(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4590_ (.A1(_0713_),
    .A2(_0692_),
    .A3(_0783_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4591_ (.A1(_0784_),
    .A2(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4592_ (.A1(_0712_),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4593_ (.I0(\dspArea_regP[12] ),
    .I1(_0787_),
    .S(_0441_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4594_ (.A1(_0355_),
    .A2(_0788_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4595_ (.A1(_2982_),
    .A2(_2988_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _4596_ (.A1(net125),
    .A2(_2987_),
    .A3(_0246_),
    .A4(_0789_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4597_ (.A1(_0248_),
    .A2(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4598_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4599_ (.A1(_0711_),
    .A2(_0786_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4600_ (.A1(_0785_),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4601_ (.A1(_0720_),
    .A2(_0782_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4602_ (.A1(_0720_),
    .A2(_0782_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4603_ (.A1(_0716_),
    .A2(_0795_),
    .A3(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4604_ (.A1(_0227_),
    .A2(_3007_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4605_ (.A1(_0644_),
    .A2(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4606_ (.A1(_0728_),
    .A2(_0741_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4607_ (.A1(_0724_),
    .A2(_0742_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4608_ (.A1(_0800_),
    .A2(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4609_ (.A1(_0799_),
    .A2(_0802_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4610_ (.I(_0739_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4611_ (.A1(_0736_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4612_ (.A1(_0731_),
    .A2(_0740_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4613_ (.A1(_0805_),
    .A2(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4614_ (.I(_0755_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4615_ (.A1(_0750_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4616_ (.A1(_0744_),
    .A2(_0745_),
    .B(_0756_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4617_ (.A1(_0809_),
    .A2(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4618_ (.A1(_0232_),
    .A2(_3000_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4619_ (.A1(_0222_),
    .A2(_3012_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4620_ (.A1(_0798_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4621_ (.A1(_0812_),
    .A2(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4622_ (.A1(_0217_),
    .A2(_3016_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4623_ (.A1(_0209_),
    .A2(_3019_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4624_ (.A1(_0205_),
    .A2(_3024_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4625_ (.A1(_0817_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4626_ (.A1(_0816_),
    .A2(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4627_ (.A1(_0211_),
    .A2(_3020_),
    .A3(_0637_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4628_ (.A1(_0218_),
    .A2(_3012_),
    .A3(_0735_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4629_ (.A1(_0821_),
    .A2(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4630_ (.A1(_0820_),
    .A2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4631_ (.A1(_0815_),
    .A2(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4632_ (.A1(_0811_),
    .A2(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4633_ (.A1(_0807_),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4634_ (.A1(_0197_),
    .A2(_3034_),
    .A3(_0657_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4635_ (.A1(_0751_),
    .A2(_0754_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4636_ (.A1(_0828_),
    .A2(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4637_ (.A1(_0758_),
    .A2(_0760_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4638_ (.A1(_0182_),
    .A2(_0177_),
    .A3(_3045_),
    .A4(_3041_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4639_ (.I(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4640_ (.A1(_0759_),
    .A2(_0831_),
    .B(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4641_ (.A1(_0200_),
    .A2(_3029_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4642_ (.A1(_0195_),
    .A2(_3032_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4643_ (.A1(_0192_),
    .A2(_3036_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4644_ (.A1(_0836_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4645_ (.A1(_0835_),
    .A2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4646_ (.A1(_0834_),
    .A2(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4647_ (.A1(_0830_),
    .A2(_0840_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4648_ (.A1(_0188_),
    .A2(_3041_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4649_ (.A1(_0181_),
    .A2(_3044_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4650_ (.A1(_0177_),
    .A2(_3048_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4651_ (.A1(_0843_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4652_ (.A1(_0842_),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4653_ (.I(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4654_ (.A1(_0173_),
    .A2(_3053_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4655_ (.A1(_0167_),
    .A2(_3057_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4656_ (.A1(\dspArea_regP[13] ),
    .A2(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4657_ (.A1(_0848_),
    .A2(_0850_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4658_ (.A1(\dspArea_regP[12] ),
    .A2(_0764_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4659_ (.A1(_0763_),
    .A2(_0765_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4660_ (.A1(_0847_),
    .A2(_0851_),
    .A3(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4661_ (.A1(_0766_),
    .A2(_0768_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4662_ (.A1(_0766_),
    .A2(_0768_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4663_ (.A1(_0762_),
    .A2(_0855_),
    .B(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4664_ (.A1(_0854_),
    .A2(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4665_ (.A1(_0841_),
    .A2(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4666_ (.A1(_0769_),
    .A2(_0772_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4667_ (.A1(_0757_),
    .A2(_0773_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4668_ (.A1(_0860_),
    .A2(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4669_ (.A1(_0827_),
    .A2(_0859_),
    .A3(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4670_ (.A1(_0775_),
    .A2(_0776_),
    .A3(_0774_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4671_ (.A1(_0775_),
    .A2(_0776_),
    .B(_0774_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4672_ (.A1(_0743_),
    .A2(_0864_),
    .B(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4673_ (.A1(_0863_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4674_ (.A1(_0803_),
    .A2(_0867_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4675_ (.A1(_0778_),
    .A2(_0781_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4676_ (.A1(_0869_),
    .A2(_0796_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4677_ (.A1(_0868_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4678_ (.A1(_0797_),
    .A2(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4679_ (.A1(_0794_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4680_ (.I(_0250_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4681_ (.A1(\dspArea_regP[13] ),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4682_ (.A1(_0792_),
    .A2(_0873_),
    .B(_0875_),
    .C(_0157_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4683_ (.A1(_0868_),
    .A2(_0870_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4684_ (.A1(_0644_),
    .A2(_0798_),
    .A3(_0802_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4685_ (.A1(_0811_),
    .A2(_0825_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4686_ (.A1(_0807_),
    .A2(_0826_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4687_ (.A1(_0878_),
    .A2(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4688_ (.A1(_0226_),
    .A2(_3011_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4689_ (.A1(_0729_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4690_ (.A1(_0234_),
    .A2(_3001_),
    .A3(_0814_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4691_ (.A1(_0882_),
    .A2(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4692_ (.A1(_0238_),
    .A2(_3002_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4693_ (.A1(_0884_),
    .A2(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4694_ (.A1(_0880_),
    .A2(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4695_ (.I(_0823_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4696_ (.A1(_0820_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4697_ (.A1(_0815_),
    .A2(_0824_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4698_ (.A1(_0889_),
    .A2(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4699_ (.I(_0839_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4700_ (.A1(_0834_),
    .A2(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4701_ (.A1(_0830_),
    .A2(_0840_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4702_ (.A1(_0893_),
    .A2(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4703_ (.A1(_0232_),
    .A2(_3008_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4704_ (.A1(_0222_),
    .A2(_3015_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4705_ (.A1(_0881_),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4706_ (.A1(_0896_),
    .A2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4707_ (.A1(_0216_),
    .A2(_3019_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4708_ (.A1(_0209_),
    .A2(_3024_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4709_ (.A1(_0205_),
    .A2(_3028_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4710_ (.A1(_0901_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4711_ (.A1(_0900_),
    .A2(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4712_ (.A1(_0211_),
    .A2(_3025_),
    .A3(_0734_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4713_ (.A1(_0217_),
    .A2(_3016_),
    .A3(_0819_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4714_ (.A1(_0905_),
    .A2(_0906_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4715_ (.A1(_0904_),
    .A2(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4716_ (.A1(_0899_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4717_ (.A1(_0895_),
    .A2(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4718_ (.A1(_0891_),
    .A2(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4719_ (.A1(_0197_),
    .A2(_3038_),
    .A3(_0753_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4720_ (.A1(_0835_),
    .A2(_0838_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4721_ (.A1(_0912_),
    .A2(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4722_ (.A1(_0183_),
    .A2(_3049_),
    .A3(_0760_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4723_ (.A1(_0189_),
    .A2(_3041_),
    .A3(_0845_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4724_ (.A1(_0404_),
    .A2(_3033_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4725_ (.A1(_0364_),
    .A2(_3036_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4726_ (.A1(_0192_),
    .A2(_3040_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4727_ (.A1(_0918_),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4728_ (.A1(_0917_),
    .A2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4729_ (.A1(_0915_),
    .A2(_0916_),
    .A3(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4730_ (.A1(_0915_),
    .A2(_0916_),
    .B(_0921_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4731_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4732_ (.A1(_0914_),
    .A2(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4733_ (.A1(_0187_),
    .A2(_3045_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4734_ (.A1(_0180_),
    .A2(_3048_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4735_ (.A1(_0176_),
    .A2(_3052_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4736_ (.A1(_0927_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4737_ (.A1(_0926_),
    .A2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4738_ (.I(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4739_ (.A1(_0173_),
    .A2(_3057_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4740_ (.A1(_0167_),
    .A2(_3060_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4741_ (.A1(\dspArea_regP[14] ),
    .A2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4742_ (.A1(_0932_),
    .A2(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4743_ (.A1(\dspArea_regP[13] ),
    .A2(_0849_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4744_ (.A1(_0848_),
    .A2(_0850_),
    .B(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4745_ (.A1(_0931_),
    .A2(_0935_),
    .A3(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4746_ (.A1(_0851_),
    .A2(_0853_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4747_ (.A1(_0851_),
    .A2(_0853_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4748_ (.A1(_0847_),
    .A2(_0939_),
    .B(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4749_ (.A1(_0938_),
    .A2(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4750_ (.A1(_0925_),
    .A2(_0942_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4751_ (.A1(_0854_),
    .A2(_0857_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4752_ (.A1(_0841_),
    .A2(_0858_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4753_ (.A1(_0944_),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4754_ (.A1(_0911_),
    .A2(_0943_),
    .A3(_0946_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4755_ (.A1(_0860_),
    .A2(_0861_),
    .A3(_0859_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4756_ (.A1(_0860_),
    .A2(_0861_),
    .B(_0859_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4757_ (.A1(_0827_),
    .A2(_0948_),
    .B(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4758_ (.A1(_0887_),
    .A2(_0947_),
    .A3(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4759_ (.A1(_0863_),
    .A2(_0866_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4760_ (.A1(_0803_),
    .A2(_0867_),
    .B(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4761_ (.A1(_0877_),
    .A2(_0951_),
    .A3(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4762_ (.A1(_0876_),
    .A2(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4763_ (.A1(_0786_),
    .A2(_0872_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4764_ (.A1(_0797_),
    .A2(_0785_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4765_ (.A1(_0871_),
    .A2(_0957_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4766_ (.A1(_0712_),
    .A2(_0956_),
    .B(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4767_ (.A1(_0955_),
    .A2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4768_ (.A1(\dspArea_regP[14] ),
    .A2(_0299_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4769_ (.A1(_0299_),
    .A2(_0960_),
    .B(_0961_),
    .C(_0157_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4770_ (.A1(\dspArea_regP[15] ),
    .A2(_0259_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4771_ (.A1(_0951_),
    .A2(_0953_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4772_ (.A1(_0951_),
    .A2(_0953_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4773_ (.A1(_0877_),
    .A2(_0963_),
    .B(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4774_ (.A1(_0880_),
    .A2(_0886_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4775_ (.A1(_0884_),
    .A2(_0885_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4776_ (.A1(_0895_),
    .A2(_0909_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4777_ (.A1(_0891_),
    .A2(_0910_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4778_ (.A1(_0968_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4779_ (.A1(_0228_),
    .A2(_3017_),
    .A3(_0813_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4780_ (.I(_0233_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4781_ (.A1(_0972_),
    .A2(_3009_),
    .A3(_0898_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4782_ (.A1(_0236_),
    .A2(_3009_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4783_ (.A1(_0971_),
    .A2(_0973_),
    .A3(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4784_ (.A1(_0971_),
    .A2(_0973_),
    .B(_0974_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4785_ (.A1(_0975_),
    .A2(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4786_ (.A1(_0241_),
    .A2(_3001_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4787_ (.A1(_0977_),
    .A2(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4788_ (.I(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4789_ (.A1(_0967_),
    .A2(_0970_),
    .A3(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4790_ (.A1(_0904_),
    .A2(_0907_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4791_ (.A1(_0899_),
    .A2(_0908_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4792_ (.A1(_0915_),
    .A2(_0916_),
    .A3(_0921_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4793_ (.A1(_0914_),
    .A2(_0984_),
    .B(_0923_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4794_ (.A1(\dspArea_regB[13] ),
    .A2(_3011_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4795_ (.A1(_0225_),
    .A2(_3015_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4796_ (.A1(_0221_),
    .A2(_3019_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4797_ (.A1(_0987_),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4798_ (.A1(_0986_),
    .A2(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4799_ (.A1(_0216_),
    .A2(_3024_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4800_ (.A1(_0209_),
    .A2(_3028_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4801_ (.A1(_0205_),
    .A2(_3032_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4802_ (.A1(_0992_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4803_ (.A1(_0991_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4804_ (.A1(_0211_),
    .A2(_3029_),
    .A3(_0818_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4805_ (.A1(_0218_),
    .A2(_3020_),
    .A3(_0903_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4806_ (.A1(_0996_),
    .A2(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4807_ (.A1(_0990_),
    .A2(_0995_),
    .A3(_0998_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4808_ (.A1(_0985_),
    .A2(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4809_ (.A1(_0982_),
    .A2(_0983_),
    .A3(_1000_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4810_ (.A1(_0982_),
    .A2(_0983_),
    .B(_1000_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4811_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4812_ (.A1(_0198_),
    .A2(_3042_),
    .A3(_0837_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4813_ (.A1(_0203_),
    .A2(_3034_),
    .A3(_0920_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4814_ (.A1(_1004_),
    .A2(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4815_ (.A1(_0184_),
    .A2(_3054_),
    .A3(_0844_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4816_ (.A1(_0190_),
    .A2(_3046_),
    .A3(_0929_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4817_ (.A1(_0201_),
    .A2(_3038_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4818_ (.A1(_0196_),
    .A2(_3040_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4819_ (.A1(_0406_),
    .A2(_3044_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4820_ (.A1(_1010_),
    .A2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4821_ (.A1(_1009_),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4822_ (.A1(_1007_),
    .A2(_1008_),
    .A3(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4823_ (.A1(_1007_),
    .A2(_1008_),
    .B(_1013_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4824_ (.A1(_1014_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4825_ (.A1(_1006_),
    .A2(_1016_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4826_ (.A1(_0186_),
    .A2(_3048_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4827_ (.A1(_0180_),
    .A2(_3052_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4828_ (.A1(_0176_),
    .A2(_3056_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4829_ (.A1(_1019_),
    .A2(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4830_ (.A1(_1018_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4831_ (.I(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4832_ (.A1(_0173_),
    .A2(_3061_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4833_ (.A1(_0529_),
    .A2(_3064_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4834_ (.A1(\dspArea_regP[15] ),
    .A2(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4835_ (.A1(_1024_),
    .A2(_1026_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4836_ (.A1(\dspArea_regP[14] ),
    .A2(_0933_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4837_ (.A1(_0932_),
    .A2(_0934_),
    .B(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4838_ (.A1(_1023_),
    .A2(_1027_),
    .A3(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4839_ (.A1(_0935_),
    .A2(_0937_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4840_ (.A1(_0935_),
    .A2(_0937_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4841_ (.A1(_0931_),
    .A2(_1031_),
    .B(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4842_ (.A1(_1030_),
    .A2(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4843_ (.A1(_1017_),
    .A2(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4844_ (.A1(_0938_),
    .A2(_0941_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4845_ (.A1(_0925_),
    .A2(_0942_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4846_ (.A1(_1036_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4847_ (.A1(_1003_),
    .A2(_1035_),
    .A3(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4848_ (.A1(_0944_),
    .A2(_0945_),
    .A3(_0943_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4849_ (.A1(_0944_),
    .A2(_0945_),
    .B(_0943_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4850_ (.A1(_0911_),
    .A2(_1040_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4851_ (.A1(_0981_),
    .A2(_1039_),
    .A3(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4852_ (.A1(_0947_),
    .A2(_0950_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4853_ (.A1(_0947_),
    .A2(_0950_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4854_ (.A1(_0887_),
    .A2(_1044_),
    .B(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4855_ (.A1(_0966_),
    .A2(_1043_),
    .A3(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4856_ (.A1(_0965_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4857_ (.A1(_0876_),
    .A2(_0954_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4858_ (.I(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4859_ (.A1(_0955_),
    .A2(_0959_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4860_ (.A1(_1050_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4861_ (.A1(_1048_),
    .A2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4862_ (.A1(_0792_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4863_ (.A1(_3173_),
    .A2(_0962_),
    .A3(_1054_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4864_ (.I(_1047_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4865_ (.A1(_0965_),
    .A2(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4866_ (.A1(_0955_),
    .A2(_1048_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4867_ (.A1(_0871_),
    .A2(_0957_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4868_ (.A1(_0965_),
    .A2(_1055_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4869_ (.I(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4870_ (.A1(_1049_),
    .A2(_1056_),
    .B1(_1057_),
    .B2(_1058_),
    .C(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4871_ (.A1(_0555_),
    .A2(_0559_),
    .B(_0618_),
    .C(_0694_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4872_ (.A1(_0708_),
    .A2(_0709_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4873_ (.A1(_0786_),
    .A2(_0872_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4874_ (.A1(_1062_),
    .A2(_1063_),
    .B(_1064_),
    .C(_1057_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4875_ (.A1(_1061_),
    .A2(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4876_ (.A1(_0970_),
    .A2(_0980_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4877_ (.A1(_0970_),
    .A2(_0980_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4878_ (.A1(_0967_),
    .A2(_1068_),
    .A3(_1067_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4879_ (.A1(_1067_),
    .A2(_1069_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4880_ (.A1(_0242_),
    .A2(_3002_),
    .A3(_0977_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4881_ (.A1(_0976_),
    .A2(_1071_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4882_ (.I(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4883_ (.A1(_0914_),
    .A2(_0924_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4884_ (.A1(_0923_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4885_ (.A1(_1075_),
    .A2(_0999_),
    .B(_1002_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4886_ (.A1(_0227_),
    .A2(_3021_),
    .A3(_0897_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4887_ (.A1(_0233_),
    .A2(_3013_),
    .A3(_0989_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4888_ (.A1(_0236_),
    .A2(_3013_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4889_ (.A1(_1077_),
    .A2(_1078_),
    .A3(_1079_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4890_ (.A1(_1077_),
    .A2(_1078_),
    .B(_1079_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4891_ (.A1(_1080_),
    .A2(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4892_ (.A1(_0240_),
    .A2(_3009_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4893_ (.A1(_1082_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4894_ (.A1(_1076_),
    .A2(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4895_ (.A1(_1073_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4896_ (.I(_0998_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4897_ (.A1(_0995_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4898_ (.A1(_0995_),
    .A2(_0998_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4899_ (.A1(_0990_),
    .A2(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4900_ (.A1(_1007_),
    .A2(_1008_),
    .A3(_1013_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4901_ (.A1(_1006_),
    .A2(_1091_),
    .B(_1015_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4902_ (.A1(_0231_),
    .A2(_3016_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4903_ (.A1(_0226_),
    .A2(_3019_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4904_ (.A1(_0221_),
    .A2(_3024_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4905_ (.A1(_1094_),
    .A2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4906_ (.A1(_1093_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4907_ (.A1(_0217_),
    .A2(_3029_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4908_ (.A1(_0210_),
    .A2(_3032_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4909_ (.A1(_0206_),
    .A2(_3036_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4910_ (.A1(_1099_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4911_ (.A1(_1098_),
    .A2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4912_ (.A1(_0212_),
    .A2(_3033_),
    .A3(_0902_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4913_ (.A1(_0634_),
    .A2(_3025_),
    .A3(_0994_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4914_ (.A1(_1103_),
    .A2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4915_ (.A1(_1097_),
    .A2(_1102_),
    .A3(_1105_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4916_ (.A1(_1092_),
    .A2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4917_ (.A1(_1088_),
    .A2(_1090_),
    .A3(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4918_ (.A1(_1088_),
    .A2(_1090_),
    .B(_1107_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4919_ (.A1(_1108_),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4920_ (.A1(_0197_),
    .A2(_3046_),
    .A3(_0919_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4921_ (.A1(_0202_),
    .A2(_3038_),
    .A3(_1012_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4922_ (.A1(_1111_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4923_ (.A1(_0183_),
    .A2(_3058_),
    .A3(_0928_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4924_ (.A1(_0189_),
    .A2(_3050_),
    .A3(_1021_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4925_ (.A1(_0404_),
    .A2(_3041_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4926_ (.A1(_0364_),
    .A2(_3044_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4927_ (.A1(_0406_),
    .A2(_3048_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4928_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4929_ (.A1(_1116_),
    .A2(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4930_ (.A1(_1114_),
    .A2(_1115_),
    .A3(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4931_ (.A1(_1114_),
    .A2(_1115_),
    .B(_1120_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4932_ (.A1(_1121_),
    .A2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4933_ (.A1(_1113_),
    .A2(_1123_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4934_ (.A1(_0186_),
    .A2(_3053_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4935_ (.A1(_0180_),
    .A2(_3056_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4936_ (.A1(\dspArea_regB[2] ),
    .A2(_3060_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4937_ (.A1(_1126_),
    .A2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4938_ (.A1(_1125_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4939_ (.I(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4940_ (.A1(_0172_),
    .A2(_3065_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4941_ (.A1(_0529_),
    .A2(_3068_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4942_ (.A1(\dspArea_regP[16] ),
    .A2(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4943_ (.A1(_1131_),
    .A2(_1133_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4944_ (.A1(\dspArea_regP[15] ),
    .A2(_1025_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4945_ (.A1(_1024_),
    .A2(_1026_),
    .B(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4946_ (.A1(_1130_),
    .A2(_1134_),
    .A3(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4947_ (.A1(_1027_),
    .A2(_1029_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4948_ (.A1(_1027_),
    .A2(_1029_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4949_ (.A1(_1023_),
    .A2(_1138_),
    .B(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4950_ (.A1(_1137_),
    .A2(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4951_ (.A1(_1124_),
    .A2(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4952_ (.A1(_1030_),
    .A2(_1033_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4953_ (.A1(_1017_),
    .A2(_1034_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4954_ (.A1(_1143_),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4955_ (.A1(_1110_),
    .A2(_1142_),
    .A3(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4956_ (.A1(_1036_),
    .A2(_1037_),
    .A3(_1035_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4957_ (.A1(_1036_),
    .A2(_1037_),
    .B(_1035_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4958_ (.A1(_1003_),
    .A2(_1147_),
    .B(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _4959_ (.A1(_1086_),
    .A2(_1146_),
    .A3(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4960_ (.A1(_1039_),
    .A2(_1042_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4961_ (.A1(_1039_),
    .A2(_1042_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4962_ (.A1(_0981_),
    .A2(_1151_),
    .B(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4963_ (.A1(_1150_),
    .A2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4964_ (.A1(_1070_),
    .A2(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4965_ (.A1(_1043_),
    .A2(_1046_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4966_ (.A1(_1043_),
    .A2(_1046_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4967_ (.A1(_0880_),
    .A2(_0886_),
    .A3(_1156_),
    .B(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4968_ (.A1(_1155_),
    .A2(_1158_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4969_ (.A1(_1066_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4970_ (.I0(\dspArea_regP[16] ),
    .I1(_1160_),
    .S(_0441_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4971_ (.A1(_0355_),
    .A2(_1161_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4972_ (.A1(\dspArea_regP[17] ),
    .A2(_0259_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4973_ (.A1(_1150_),
    .A2(_1153_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4974_ (.A1(_1070_),
    .A2(_1154_),
    .B(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4975_ (.A1(_1076_),
    .A2(_1084_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4976_ (.A1(_1073_),
    .A2(_1085_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4977_ (.A1(_1165_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4978_ (.A1(_0244_),
    .A2(_3009_),
    .A3(_1082_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4979_ (.A1(_1081_),
    .A2(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4980_ (.A1(_1006_),
    .A2(_1016_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4981_ (.A1(_1015_),
    .A2(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4982_ (.A1(_1171_),
    .A2(_1106_),
    .B(_1109_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4983_ (.A1(_0229_),
    .A2(_3026_),
    .A3(_0988_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4984_ (.A1(_0972_),
    .A2(_3017_),
    .A3(_1096_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4985_ (.A1(_0237_),
    .A2(_3017_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4986_ (.A1(_1173_),
    .A2(_1174_),
    .A3(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4987_ (.A1(_1173_),
    .A2(_1174_),
    .B(_1175_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4988_ (.A1(_1176_),
    .A2(_1177_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4989_ (.A1(_0241_),
    .A2(_3013_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4990_ (.A1(_1178_),
    .A2(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4991_ (.A1(_1172_),
    .A2(_1180_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4992_ (.A1(_1169_),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4993_ (.I(_1105_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4994_ (.A1(_1102_),
    .A2(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4995_ (.A1(_1102_),
    .A2(_1105_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4996_ (.A1(_1097_),
    .A2(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4997_ (.A1(_1114_),
    .A2(_1115_),
    .A3(_1120_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4998_ (.A1(_1113_),
    .A2(_1187_),
    .B(_1122_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4999_ (.A1(_0231_),
    .A2(_3020_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5000_ (.A1(_0225_),
    .A2(_3024_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5001_ (.A1(_0221_),
    .A2(_3028_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5002_ (.A1(_1190_),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5003_ (.A1(_1189_),
    .A2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5004_ (.A1(_0216_),
    .A2(_3033_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5005_ (.A1(_0209_),
    .A2(_3036_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5006_ (.A1(_0205_),
    .A2(_3040_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5007_ (.A1(_1195_),
    .A2(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5008_ (.A1(_1194_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5009_ (.A1(_0212_),
    .A2(_3037_),
    .A3(_0993_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5010_ (.A1(_0218_),
    .A2(_3029_),
    .A3(_1101_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5011_ (.A1(_1199_),
    .A2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5012_ (.A1(_1193_),
    .A2(_1198_),
    .A3(_1201_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5013_ (.A1(_1188_),
    .A2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5014_ (.A1(_1184_),
    .A2(_1186_),
    .A3(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5015_ (.A1(_1184_),
    .A2(_1186_),
    .B(_1203_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5016_ (.A1(_1204_),
    .A2(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5017_ (.A1(_0198_),
    .A2(_3050_),
    .A3(_1011_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5018_ (.A1(_0203_),
    .A2(_3042_),
    .A3(_1119_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5019_ (.A1(_1207_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5020_ (.A1(_0184_),
    .A2(_3062_),
    .A3(_1020_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5021_ (.A1(_0190_),
    .A2(_3054_),
    .A3(_1128_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5022_ (.A1(_0201_),
    .A2(_3045_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5023_ (.A1(_0196_),
    .A2(_3049_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5024_ (.A1(_0406_),
    .A2(_3052_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5025_ (.A1(_1213_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5026_ (.A1(_1212_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5027_ (.A1(_1210_),
    .A2(_1211_),
    .A3(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5028_ (.A1(_1210_),
    .A2(_1211_),
    .B(_1216_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5029_ (.A1(_1217_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5030_ (.A1(_1209_),
    .A2(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5031_ (.A1(_0186_),
    .A2(_3057_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5032_ (.A1(_0180_),
    .A2(_3060_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5033_ (.A1(_0176_),
    .A2(_3064_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5034_ (.A1(_1222_),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5035_ (.A1(_1221_),
    .A2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5036_ (.I(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5037_ (.A1(_0173_),
    .A2(_3069_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5038_ (.A1(_0529_),
    .A2(_3074_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5039_ (.A1(\dspArea_regP[17] ),
    .A2(_1228_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5040_ (.A1(_1227_),
    .A2(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5041_ (.A1(\dspArea_regP[16] ),
    .A2(_1132_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5042_ (.A1(_1131_),
    .A2(_1133_),
    .B(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5043_ (.A1(_1226_),
    .A2(_1230_),
    .A3(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5044_ (.A1(_1134_),
    .A2(_1136_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5045_ (.A1(_1134_),
    .A2(_1136_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5046_ (.A1(_1130_),
    .A2(_1234_),
    .B(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5047_ (.A1(_1233_),
    .A2(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5048_ (.A1(_1220_),
    .A2(_1237_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5049_ (.A1(_1137_),
    .A2(_1140_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5050_ (.A1(_1124_),
    .A2(_1141_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5051_ (.A1(_1239_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5052_ (.A1(_1206_),
    .A2(_1238_),
    .A3(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5053_ (.A1(_1143_),
    .A2(_1144_),
    .A3(_1142_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5054_ (.A1(_1143_),
    .A2(_1144_),
    .B(_1142_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5055_ (.A1(_1110_),
    .A2(_1243_),
    .B(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5056_ (.A1(_1242_),
    .A2(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5057_ (.A1(_1182_),
    .A2(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5058_ (.A1(_1146_),
    .A2(_1149_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5059_ (.A1(_1146_),
    .A2(_1149_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5060_ (.A1(_1086_),
    .A2(_1248_),
    .B(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5061_ (.A1(_1167_),
    .A2(_1247_),
    .A3(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5062_ (.A1(_1164_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5063_ (.A1(_1155_),
    .A2(_1158_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5064_ (.I(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5065_ (.I(_1056_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5066_ (.A1(_0955_),
    .A2(_1048_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5067_ (.A1(_1050_),
    .A2(_1255_),
    .B1(_1256_),
    .B2(_0958_),
    .C(_1059_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5068_ (.A1(_0707_),
    .A2(_0710_),
    .B(_0956_),
    .C(_1256_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5069_ (.A1(_1257_),
    .A2(_1258_),
    .B(_1159_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5070_ (.A1(_1254_),
    .A2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5071_ (.A1(_1252_),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5072_ (.A1(_0792_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5073_ (.A1(_3173_),
    .A2(_1162_),
    .A3(_1262_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5074_ (.A1(_1172_),
    .A2(_1180_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5075_ (.I(_1169_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5076_ (.A1(_1264_),
    .A2(_1181_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5077_ (.A1(_1263_),
    .A2(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5078_ (.A1(_0242_),
    .A2(_3013_),
    .A3(_1178_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5079_ (.A1(_1177_),
    .A2(_1267_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5080_ (.I(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5081_ (.A1(_1113_),
    .A2(_1123_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5082_ (.A1(_1122_),
    .A2(_1270_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5083_ (.A1(_1271_),
    .A2(_1202_),
    .B(_1205_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5084_ (.A1(_0228_),
    .A2(_3030_),
    .A3(_1095_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5085_ (.A1(_0233_),
    .A2(_3021_),
    .A3(_1192_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5086_ (.A1(_0236_),
    .A2(_3021_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5087_ (.A1(_1273_),
    .A2(_1274_),
    .A3(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5088_ (.A1(_1273_),
    .A2(_1274_),
    .B(_1275_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5089_ (.A1(_1276_),
    .A2(_1277_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5090_ (.A1(_0240_),
    .A2(_3017_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5091_ (.A1(_1278_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5092_ (.A1(_1272_),
    .A2(_1280_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5093_ (.A1(_1269_),
    .A2(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5094_ (.I(_1201_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5095_ (.A1(_1198_),
    .A2(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5096_ (.A1(_1198_),
    .A2(_1201_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5097_ (.A1(_1193_),
    .A2(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5098_ (.A1(_1210_),
    .A2(_1211_),
    .A3(_1216_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5099_ (.A1(_1209_),
    .A2(_1287_),
    .B(_1218_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5100_ (.A1(_0231_),
    .A2(_3025_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5101_ (.A1(_0226_),
    .A2(_3028_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5102_ (.A1(_0221_),
    .A2(_3032_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5103_ (.A1(_1290_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5104_ (.A1(_1289_),
    .A2(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5105_ (.A1(_0217_),
    .A2(_3037_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5106_ (.A1(_0210_),
    .A2(_3040_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5107_ (.A1(_0206_),
    .A2(_3044_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5108_ (.A1(_1295_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5109_ (.A1(_1294_),
    .A2(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5110_ (.A1(_0213_),
    .A2(_3041_),
    .A3(_1100_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5111_ (.A1(_0634_),
    .A2(_3034_),
    .A3(_1197_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5112_ (.A1(_1299_),
    .A2(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5113_ (.A1(_1293_),
    .A2(_1298_),
    .A3(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5114_ (.A1(_1288_),
    .A2(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5115_ (.A1(_1284_),
    .A2(_1286_),
    .A3(_1303_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5116_ (.A1(_1284_),
    .A2(_1286_),
    .B(_1303_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5117_ (.A1(_1304_),
    .A2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5118_ (.A1(_0197_),
    .A2(_3053_),
    .A3(_1118_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5119_ (.A1(_0202_),
    .A2(_3046_),
    .A3(_1215_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5120_ (.A1(_1307_),
    .A2(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5121_ (.A1(_0183_),
    .A2(_3065_),
    .A3(_1127_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5122_ (.A1(_0189_),
    .A2(_3058_),
    .A3(_1224_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5123_ (.A1(_0404_),
    .A2(_3049_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5124_ (.A1(_0364_),
    .A2(_3052_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5125_ (.A1(_0406_),
    .A2(_3056_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5126_ (.A1(_1313_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5127_ (.A1(_1312_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5128_ (.A1(_1310_),
    .A2(_1311_),
    .A3(_1316_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5129_ (.A1(_1310_),
    .A2(_1311_),
    .B(_1316_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5130_ (.A1(_1317_),
    .A2(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5131_ (.A1(_1309_),
    .A2(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5132_ (.A1(_0186_),
    .A2(_3061_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5133_ (.A1(_0180_),
    .A2(_3064_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5134_ (.A1(_0176_),
    .A2(_3068_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5135_ (.A1(_1322_),
    .A2(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5136_ (.A1(_1321_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5137_ (.I(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5138_ (.A1(_0173_),
    .A2(_3075_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5139_ (.A1(_0529_),
    .A2(_3079_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5140_ (.A1(\dspArea_regP[18] ),
    .A2(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5141_ (.A1(_1327_),
    .A2(_1329_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5142_ (.A1(\dspArea_regP[17] ),
    .A2(_1228_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5143_ (.A1(_1227_),
    .A2(_1229_),
    .B(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5144_ (.A1(_1326_),
    .A2(_1330_),
    .A3(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5145_ (.A1(_1230_),
    .A2(_1232_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5146_ (.A1(_1230_),
    .A2(_1232_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5147_ (.A1(_1226_),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5148_ (.A1(_1333_),
    .A2(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5149_ (.A1(_1320_),
    .A2(_1337_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5150_ (.A1(_1233_),
    .A2(_1236_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5151_ (.A1(_1220_),
    .A2(_1237_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5152_ (.A1(_1339_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5153_ (.A1(_1306_),
    .A2(_1338_),
    .A3(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5154_ (.A1(_1239_),
    .A2(_1240_),
    .A3(_1238_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5155_ (.A1(_1239_),
    .A2(_1240_),
    .B(_1238_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5156_ (.A1(_1206_),
    .A2(_1343_),
    .B(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5157_ (.A1(_1282_),
    .A2(_1342_),
    .A3(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5158_ (.A1(_1242_),
    .A2(_1245_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5159_ (.A1(_1182_),
    .A2(_1246_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5160_ (.A1(_1347_),
    .A2(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5161_ (.A1(_1266_),
    .A2(_1346_),
    .A3(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5162_ (.A1(_1247_),
    .A2(_1250_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5163_ (.A1(_1247_),
    .A2(_1250_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5164_ (.A1(_1167_),
    .A2(_1351_),
    .B(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5165_ (.A1(_1350_),
    .A2(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5166_ (.A1(_1159_),
    .A2(_1252_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5167_ (.A1(_1070_),
    .A2(_1154_),
    .B(_1251_),
    .C(_1163_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5168_ (.A1(_1155_),
    .A2(_1158_),
    .A3(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5169_ (.A1(_1167_),
    .A2(_1351_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5170_ (.A1(_1167_),
    .A2(_1351_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5171_ (.A1(_1164_),
    .A2(_1358_),
    .A3(_1359_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5172_ (.A1(_1066_),
    .A2(_1355_),
    .B(_1357_),
    .C(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5173_ (.A1(_1354_),
    .A2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5174_ (.I0(\dspArea_regP[18] ),
    .I1(_1362_),
    .S(_0441_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5175_ (.A1(_0355_),
    .A2(_1363_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5176_ (.A1(_1347_),
    .A2(_1348_),
    .A3(_1346_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5177_ (.A1(_1347_),
    .A2(_1348_),
    .B(_1346_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5178_ (.A1(_1266_),
    .A2(_1364_),
    .B(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5179_ (.A1(_1272_),
    .A2(_1280_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5180_ (.A1(_1269_),
    .A2(_1281_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5181_ (.A1(_1367_),
    .A2(_1368_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5182_ (.A1(_0243_),
    .A2(_3017_),
    .A3(_1278_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5183_ (.A1(_1277_),
    .A2(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5184_ (.A1(_1209_),
    .A2(_1219_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5185_ (.A1(_1218_),
    .A2(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5186_ (.A1(_1373_),
    .A2(_1302_),
    .B(_1305_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5187_ (.A1(_0228_),
    .A2(_3034_),
    .A3(_1191_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5188_ (.A1(_0233_),
    .A2(_3026_),
    .A3(_1292_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5189_ (.A1(_0236_),
    .A2(_3026_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5190_ (.A1(_1375_),
    .A2(_1376_),
    .A3(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5191_ (.A1(_1375_),
    .A2(_1376_),
    .B(_1377_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5192_ (.A1(_1378_),
    .A2(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5193_ (.A1(_0241_),
    .A2(_3021_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5194_ (.A1(_1380_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5195_ (.A1(_1374_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5196_ (.A1(_1371_),
    .A2(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5197_ (.I(_1301_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5198_ (.A1(_1298_),
    .A2(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5199_ (.A1(_1298_),
    .A2(_1301_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5200_ (.A1(_1293_),
    .A2(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5201_ (.A1(_1310_),
    .A2(_1311_),
    .A3(_1316_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5202_ (.A1(_1309_),
    .A2(_1389_),
    .B(_1318_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5203_ (.A1(_0231_),
    .A2(_3029_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5204_ (.A1(_0225_),
    .A2(_3032_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5205_ (.A1(_0221_),
    .A2(_3036_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5206_ (.A1(_1392_),
    .A2(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5207_ (.A1(_1391_),
    .A2(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5208_ (.A1(_0216_),
    .A2(_3040_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5209_ (.A1(_0209_),
    .A2(_3044_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5210_ (.A1(_0205_),
    .A2(_3048_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5211_ (.A1(_1397_),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5212_ (.A1(_1396_),
    .A2(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5213_ (.A1(_0212_),
    .A2(_3045_),
    .A3(_1196_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5214_ (.A1(_0218_),
    .A2(_3037_),
    .A3(_1297_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5215_ (.A1(_1401_),
    .A2(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5216_ (.A1(_1395_),
    .A2(_1400_),
    .A3(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5217_ (.A1(_1390_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5218_ (.A1(_1386_),
    .A2(_1388_),
    .A3(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5219_ (.A1(_1386_),
    .A2(_1388_),
    .B(_1405_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5220_ (.A1(_1406_),
    .A2(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5221_ (.A1(_0196_),
    .A2(_3057_),
    .A3(_1214_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5222_ (.A1(_0201_),
    .A2(_3049_),
    .A3(_1315_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5223_ (.A1(_1409_),
    .A2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5224_ (.A1(_0182_),
    .A2(_3069_),
    .A3(_1223_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5225_ (.A1(_0187_),
    .A2(_3061_),
    .A3(_1324_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5226_ (.A1(_0200_),
    .A2(_3053_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5227_ (.A1(_0195_),
    .A2(_3056_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5228_ (.A1(_0192_),
    .A2(_3060_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5229_ (.A1(_1415_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5230_ (.A1(_1414_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5231_ (.A1(_1412_),
    .A2(_1413_),
    .A3(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5232_ (.A1(_1412_),
    .A2(_1413_),
    .B(_1418_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5233_ (.A1(_1419_),
    .A2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5234_ (.A1(_1411_),
    .A2(_1421_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5235_ (.A1(_0186_),
    .A2(_3065_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5236_ (.A1(_0180_),
    .A2(_3068_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5237_ (.A1(\dspArea_regB[2] ),
    .A2(_3074_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5238_ (.A1(_1424_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5239_ (.A1(_1423_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5240_ (.I(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5241_ (.A1(_0172_),
    .A2(_3080_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5242_ (.A1(_0529_),
    .A2(_3084_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5243_ (.A1(\dspArea_regP[19] ),
    .A2(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5244_ (.A1(_1429_),
    .A2(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5245_ (.A1(\dspArea_regP[18] ),
    .A2(_1328_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5246_ (.A1(_1327_),
    .A2(_1329_),
    .B(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5247_ (.A1(_1428_),
    .A2(_1432_),
    .A3(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5248_ (.A1(_1330_),
    .A2(_1332_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5249_ (.A1(_1330_),
    .A2(_1332_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5250_ (.A1(_1326_),
    .A2(_1436_),
    .B(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5251_ (.A1(_1422_),
    .A2(_1435_),
    .A3(_1438_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5252_ (.A1(_1333_),
    .A2(_1336_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5253_ (.A1(_1320_),
    .A2(_1337_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5254_ (.A1(_1440_),
    .A2(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5255_ (.A1(_1408_),
    .A2(_1439_),
    .A3(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5256_ (.A1(_1339_),
    .A2(_1340_),
    .A3(_1338_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5257_ (.A1(_1339_),
    .A2(_1340_),
    .B(_1338_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5258_ (.A1(_1306_),
    .A2(_1444_),
    .B(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5259_ (.A1(_1443_),
    .A2(_1446_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5260_ (.A1(_1384_),
    .A2(_1447_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5261_ (.A1(_1342_),
    .A2(_1345_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5262_ (.A1(_1342_),
    .A2(_1345_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5263_ (.A1(_1282_),
    .A2(_1449_),
    .B(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5264_ (.A1(_1448_),
    .A2(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5265_ (.A1(_1369_),
    .A2(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5266_ (.A1(_1366_),
    .A2(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5267_ (.A1(_1350_),
    .A2(_1353_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5268_ (.A1(_1350_),
    .A2(_1353_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5269_ (.A1(_1456_),
    .A2(_1361_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5270_ (.A1(_1455_),
    .A2(_1457_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5271_ (.A1(_1454_),
    .A2(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5272_ (.A1(\dspArea_regP[19] ),
    .A2(_0874_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5273_ (.I(_3109_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5274_ (.A1(_0792_),
    .A2(_1459_),
    .B(_1460_),
    .C(_1461_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5275_ (.A1(_1374_),
    .A2(_1382_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5276_ (.I(_1371_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5277_ (.A1(_1463_),
    .A2(_1383_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5278_ (.A1(_1462_),
    .A2(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5279_ (.A1(_0243_),
    .A2(_3021_),
    .A3(_1380_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5280_ (.A1(_1379_),
    .A2(_1466_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5281_ (.I(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5282_ (.A1(_1309_),
    .A2(_1319_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5283_ (.A1(_1318_),
    .A2(_1469_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5284_ (.A1(_1470_),
    .A2(_1404_),
    .B(_1407_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5285_ (.A1(_0229_),
    .A2(_3038_),
    .A3(_1291_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5286_ (.A1(_0972_),
    .A2(_3030_),
    .A3(_1394_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5287_ (.A1(_0236_),
    .A2(_3030_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5288_ (.A1(_1472_),
    .A2(_1473_),
    .A3(_1474_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5289_ (.A1(_1472_),
    .A2(_1473_),
    .B(_1474_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5290_ (.A1(_1475_),
    .A2(_1476_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5291_ (.A1(_0241_),
    .A2(_3026_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5292_ (.A1(_1477_),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5293_ (.A1(_1471_),
    .A2(_1479_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5294_ (.A1(_1468_),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5295_ (.I(_1403_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5296_ (.A1(_1400_),
    .A2(_1482_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5297_ (.A1(_1400_),
    .A2(_1403_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5298_ (.A1(_1395_),
    .A2(_1484_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5299_ (.A1(_1412_),
    .A2(_1413_),
    .A3(_1418_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5300_ (.A1(_1411_),
    .A2(_1486_),
    .B(_1420_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5301_ (.A1(_0232_),
    .A2(_3033_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5302_ (.A1(_0226_),
    .A2(_3036_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5303_ (.A1(_0222_),
    .A2(_3040_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5304_ (.A1(_1489_),
    .A2(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5305_ (.A1(_1488_),
    .A2(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5306_ (.A1(_0218_),
    .A2(_3045_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5307_ (.A1(_0210_),
    .A2(_3048_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5308_ (.A1(_0206_),
    .A2(_3052_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5309_ (.A1(_1494_),
    .A2(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5310_ (.A1(_1493_),
    .A2(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5311_ (.A1(_0213_),
    .A2(_3050_),
    .A3(_1296_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5312_ (.A1(_0219_),
    .A2(_3042_),
    .A3(_1399_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5313_ (.A1(_1498_),
    .A2(_1499_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5314_ (.A1(_1492_),
    .A2(_1497_),
    .A3(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5315_ (.A1(_1487_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5316_ (.A1(_1483_),
    .A2(_1485_),
    .A3(_1502_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5317_ (.A1(_1483_),
    .A2(_1485_),
    .B(_1502_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5318_ (.A1(_1503_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5319_ (.A1(_0198_),
    .A2(_3062_),
    .A3(_1314_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5320_ (.A1(_0203_),
    .A2(_3054_),
    .A3(_1417_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5321_ (.A1(_1506_),
    .A2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5322_ (.A1(_0184_),
    .A2(_3076_),
    .A3(_1323_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5323_ (.A1(_0190_),
    .A2(_3066_),
    .A3(_1426_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5324_ (.A1(_0201_),
    .A2(_3057_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5325_ (.A1(_0196_),
    .A2(_3061_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5326_ (.A1(_0406_),
    .A2(_3065_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5327_ (.A1(_1512_),
    .A2(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5328_ (.A1(_1511_),
    .A2(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5329_ (.A1(_1509_),
    .A2(_1510_),
    .A3(_1515_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5330_ (.A1(_1509_),
    .A2(_1510_),
    .B(_1515_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5331_ (.A1(_1516_),
    .A2(_1517_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5332_ (.A1(_1508_),
    .A2(_1518_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5333_ (.A1(_0188_),
    .A2(_3069_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5334_ (.A1(_0182_),
    .A2(_3074_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5335_ (.A1(_0177_),
    .A2(_3079_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5336_ (.A1(_1521_),
    .A2(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5337_ (.A1(_1520_),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5338_ (.A1(_0172_),
    .A2(_3085_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5339_ (.A1(_0529_),
    .A2(\dspArea_regA[20] ),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5340_ (.A1(\dspArea_regP[20] ),
    .A2(_1526_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5341_ (.A1(_1525_),
    .A2(_1527_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5342_ (.A1(\dspArea_regP[19] ),
    .A2(_1430_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5343_ (.A1(_1429_),
    .A2(_1431_),
    .B(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5344_ (.A1(_1528_),
    .A2(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5345_ (.A1(_1524_),
    .A2(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5346_ (.A1(_1432_),
    .A2(_1434_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5347_ (.A1(_1432_),
    .A2(_1434_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5348_ (.A1(_1428_),
    .A2(_1533_),
    .B(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5349_ (.A1(_1532_),
    .A2(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5350_ (.A1(_1519_),
    .A2(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5351_ (.A1(_1435_),
    .A2(_1438_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5352_ (.A1(_1435_),
    .A2(_1438_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5353_ (.A1(_1422_),
    .A2(_1538_),
    .B(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5354_ (.A1(_1537_),
    .A2(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5355_ (.A1(_1505_),
    .A2(_1541_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5356_ (.A1(_1440_),
    .A2(_1441_),
    .A3(_1439_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5357_ (.A1(_1440_),
    .A2(_1441_),
    .B(_1439_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5358_ (.A1(_1408_),
    .A2(_1543_),
    .B(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5359_ (.A1(_1481_),
    .A2(_1542_),
    .A3(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5360_ (.A1(_1443_),
    .A2(_1446_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5361_ (.A1(_1384_),
    .A2(_1447_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5362_ (.A1(_1547_),
    .A2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5363_ (.A1(_1465_),
    .A2(_1546_),
    .A3(_1549_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5364_ (.A1(_1448_),
    .A2(_1451_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5365_ (.A1(_1369_),
    .A2(_1452_),
    .B(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5366_ (.A1(_1550_),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5367_ (.A1(_1550_),
    .A2(_1552_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5368_ (.A1(_1553_),
    .A2(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5369_ (.A1(_1366_),
    .A2(_1453_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5370_ (.A1(_1366_),
    .A2(_1453_),
    .B(_1350_),
    .C(_1353_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5371_ (.A1(_1556_),
    .A2(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5372_ (.A1(_1360_),
    .A2(_1357_),
    .B(_1454_),
    .C(_1354_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5373_ (.A1(_1366_),
    .A2(_1453_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5374_ (.A1(_1456_),
    .A2(_1560_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5375_ (.I(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5376_ (.A1(_1061_),
    .A2(_1065_),
    .B(_1355_),
    .C(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5377_ (.A1(_1558_),
    .A2(_1559_),
    .A3(_1563_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5378_ (.A1(_1555_),
    .A2(_1564_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5379_ (.I0(\dspArea_regP[20] ),
    .I1(_1565_),
    .S(_0441_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5380_ (.A1(_0355_),
    .A2(_1566_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5381_ (.I(\dspArea_regP[21] ),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5382_ (.A1(_1555_),
    .A2(_1564_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5383_ (.A1(_1547_),
    .A2(_1548_),
    .A3(_1546_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5384_ (.A1(_1547_),
    .A2(_1548_),
    .B(_1546_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5385_ (.A1(_1465_),
    .A2(_1569_),
    .B(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5386_ (.A1(_1471_),
    .A2(_1479_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5387_ (.A1(_1468_),
    .A2(_1480_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5388_ (.A1(_1572_),
    .A2(_1573_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5389_ (.A1(_0244_),
    .A2(_3026_),
    .A3(_1477_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5390_ (.A1(_1476_),
    .A2(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5391_ (.A1(_1411_),
    .A2(_1421_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5392_ (.A1(_1420_),
    .A2(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5393_ (.A1(_1578_),
    .A2(_1501_),
    .B(_1504_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5394_ (.A1(_0229_),
    .A2(_3042_),
    .A3(_1393_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5395_ (.A1(_0972_),
    .A2(_3034_),
    .A3(_1491_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5396_ (.A1(_0237_),
    .A2(_3034_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5397_ (.A1(_1580_),
    .A2(_1581_),
    .A3(_1582_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5398_ (.A1(_1580_),
    .A2(_1581_),
    .B(_1582_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5399_ (.A1(_1583_),
    .A2(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5400_ (.A1(_0241_),
    .A2(_3030_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5401_ (.A1(_1585_),
    .A2(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5402_ (.A1(_1579_),
    .A2(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5403_ (.A1(_1576_),
    .A2(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5404_ (.I(_1500_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5405_ (.A1(_1497_),
    .A2(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5406_ (.A1(_1497_),
    .A2(_1500_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5407_ (.A1(_1492_),
    .A2(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5408_ (.A1(_1509_),
    .A2(_1510_),
    .A3(_1515_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5409_ (.A1(_1508_),
    .A2(_1594_),
    .B(_1517_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5410_ (.A1(_0231_),
    .A2(_3037_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5411_ (.A1(_0226_),
    .A2(_3040_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5412_ (.A1(_0222_),
    .A2(_3044_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5413_ (.A1(_1597_),
    .A2(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5414_ (.A1(_1596_),
    .A2(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5415_ (.A1(_0217_),
    .A2(_3049_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5416_ (.A1(_0210_),
    .A2(_3052_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5417_ (.A1(_0206_),
    .A2(_3056_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5418_ (.A1(_1602_),
    .A2(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5419_ (.A1(_1601_),
    .A2(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5420_ (.A1(_0213_),
    .A2(_3053_),
    .A3(_1398_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5421_ (.A1(_0634_),
    .A2(_3045_),
    .A3(_1496_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5422_ (.A1(_1606_),
    .A2(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5423_ (.A1(_1600_),
    .A2(_1605_),
    .A3(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5424_ (.A1(_1595_),
    .A2(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5425_ (.A1(_1591_),
    .A2(_1593_),
    .A3(_1610_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5426_ (.A1(_1591_),
    .A2(_1593_),
    .B(_1610_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5427_ (.A1(_1611_),
    .A2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5428_ (.A1(_0197_),
    .A2(_3066_),
    .A3(_1416_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5429_ (.A1(_0202_),
    .A2(_3058_),
    .A3(_1514_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5430_ (.A1(_1614_),
    .A2(_1615_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5431_ (.A1(_0183_),
    .A2(_3081_),
    .A3(_1425_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5432_ (.A1(_0189_),
    .A2(_3070_),
    .A3(_1523_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5433_ (.A1(_0404_),
    .A2(_3061_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5434_ (.A1(_0364_),
    .A2(_3065_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5435_ (.A1(_0406_),
    .A2(_3068_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5436_ (.A1(_1620_),
    .A2(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5437_ (.A1(_1619_),
    .A2(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5438_ (.A1(_1617_),
    .A2(_1618_),
    .A3(_1623_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5439_ (.A1(_1617_),
    .A2(_1618_),
    .B(_1623_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5440_ (.A1(_1624_),
    .A2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5441_ (.A1(_1616_),
    .A2(_1626_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5442_ (.A1(_0187_),
    .A2(_3075_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5443_ (.A1(_0180_),
    .A2(_3079_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5444_ (.A1(_0176_),
    .A2(_3084_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5445_ (.A1(_1629_),
    .A2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5446_ (.A1(_1628_),
    .A2(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5447_ (.A1(_0172_),
    .A2(_3089_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5448_ (.A1(_0529_),
    .A2(\dspArea_regA[21] ),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5449_ (.A1(\dspArea_regP[21] ),
    .A2(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5450_ (.A1(_1633_),
    .A2(_1635_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5451_ (.A1(\dspArea_regP[20] ),
    .A2(_1526_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5452_ (.A1(_1525_),
    .A2(_1527_),
    .B(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5453_ (.A1(_1632_),
    .A2(_1636_),
    .A3(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5454_ (.I(_1524_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5455_ (.A1(_1528_),
    .A2(_1530_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5456_ (.A1(_1528_),
    .A2(_1530_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5457_ (.A1(_1640_),
    .A2(_1641_),
    .B(_1642_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5458_ (.A1(_1639_),
    .A2(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5459_ (.A1(_1627_),
    .A2(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5460_ (.A1(_1524_),
    .A2(_1531_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5461_ (.A1(_1524_),
    .A2(_1531_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5462_ (.A1(_1646_),
    .A2(_1647_),
    .A3(_1535_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5463_ (.A1(_1519_),
    .A2(_1536_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5464_ (.A1(_1648_),
    .A2(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5465_ (.A1(_1613_),
    .A2(_1645_),
    .A3(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5466_ (.A1(_1537_),
    .A2(_1540_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5467_ (.A1(_1505_),
    .A2(_1541_),
    .B(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5468_ (.A1(_1651_),
    .A2(_1653_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5469_ (.A1(_1589_),
    .A2(_1654_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5470_ (.A1(_1542_),
    .A2(_1545_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5471_ (.A1(_1542_),
    .A2(_1545_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5472_ (.A1(_1481_),
    .A2(_1656_),
    .B(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5473_ (.A1(_1574_),
    .A2(_1655_),
    .A3(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5474_ (.A1(_1571_),
    .A2(_1659_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5475_ (.A1(_1554_),
    .A2(_1568_),
    .A3(_1660_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5476_ (.A1(_1554_),
    .A2(_1568_),
    .B(_1660_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5477_ (.A1(_0792_),
    .A2(_1661_),
    .A3(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5478_ (.A1(_1567_),
    .A2(_0297_),
    .B(_1663_),
    .C(_1461_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5479_ (.A1(_1579_),
    .A2(_1587_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5480_ (.I(_1576_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5481_ (.A1(_1665_),
    .A2(_1588_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5482_ (.A1(_1664_),
    .A2(_1666_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5483_ (.A1(_0244_),
    .A2(_3030_),
    .A3(_1585_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5484_ (.A1(_1584_),
    .A2(_1668_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5485_ (.A1(_1508_),
    .A2(_1518_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5486_ (.A1(_1517_),
    .A2(_1670_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5487_ (.A1(_1671_),
    .A2(_1609_),
    .B(_1612_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5488_ (.A1(_0229_),
    .A2(_3046_),
    .A3(_1490_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5489_ (.A1(_0972_),
    .A2(_3038_),
    .A3(_1599_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5490_ (.A1(_0237_),
    .A2(_3038_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5491_ (.A1(_1673_),
    .A2(_1674_),
    .A3(_1675_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5492_ (.A1(_1673_),
    .A2(_1674_),
    .B(_1675_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5493_ (.A1(_1676_),
    .A2(_1677_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5494_ (.A1(_0241_),
    .A2(_3034_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5495_ (.A1(_1678_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5496_ (.A1(_1672_),
    .A2(_1680_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5497_ (.A1(_1669_),
    .A2(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5498_ (.I(_1608_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5499_ (.A1(_1605_),
    .A2(_1683_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5500_ (.A1(_1605_),
    .A2(_1608_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5501_ (.A1(_1600_),
    .A2(_1685_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5502_ (.A1(_1617_),
    .A2(_1618_),
    .A3(_1623_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5503_ (.A1(_1616_),
    .A2(_1687_),
    .B(_1625_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5504_ (.A1(_0231_),
    .A2(_3041_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5505_ (.A1(_0226_),
    .A2(_3044_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5506_ (.A1(_0221_),
    .A2(_3048_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5507_ (.A1(_1690_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5508_ (.A1(_1689_),
    .A2(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5509_ (.A1(_0216_),
    .A2(_3053_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5510_ (.A1(_0209_),
    .A2(_3056_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5511_ (.A1(_0205_),
    .A2(_3060_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5512_ (.A1(_1695_),
    .A2(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5513_ (.A1(_1694_),
    .A2(_1697_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5514_ (.A1(_0212_),
    .A2(_3057_),
    .A3(_1495_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5515_ (.A1(_0634_),
    .A2(_3049_),
    .A3(_1604_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5516_ (.A1(_1699_),
    .A2(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5517_ (.A1(_1693_),
    .A2(_1698_),
    .A3(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5518_ (.A1(_1688_),
    .A2(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5519_ (.A1(_1684_),
    .A2(_1686_),
    .A3(_1703_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5520_ (.A1(_1684_),
    .A2(_1686_),
    .B(_1703_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5521_ (.A1(_1704_),
    .A2(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5522_ (.A1(_0197_),
    .A2(_3070_),
    .A3(_1513_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5523_ (.A1(_0202_),
    .A2(_3062_),
    .A3(_1622_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5524_ (.A1(_1707_),
    .A2(_1708_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5525_ (.A1(_0183_),
    .A2(_3085_),
    .A3(_1522_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5526_ (.A1(_0189_),
    .A2(_3076_),
    .A3(_1631_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5527_ (.A1(_0404_),
    .A2(_3065_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5528_ (.A1(_0364_),
    .A2(_3069_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5529_ (.A1(_0406_),
    .A2(_3074_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5530_ (.A1(_1713_),
    .A2(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5531_ (.A1(_1712_),
    .A2(_1715_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5532_ (.A1(_1710_),
    .A2(_1711_),
    .A3(_1716_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5533_ (.A1(_1710_),
    .A2(_1711_),
    .B(_1716_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5534_ (.A1(_1717_),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5535_ (.A1(_1709_),
    .A2(_1719_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5536_ (.A1(_0186_),
    .A2(_3080_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5537_ (.A1(_0180_),
    .A2(_3084_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5538_ (.A1(\dspArea_regB[2] ),
    .A2(\dspArea_regA[20] ),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5539_ (.A1(_1722_),
    .A2(_1723_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5540_ (.A1(_1721_),
    .A2(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5541_ (.I(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5542_ (.A1(_0172_),
    .A2(_3093_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5543_ (.A1(_0529_),
    .A2(\dspArea_regA[22] ),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5544_ (.A1(\dspArea_regP[22] ),
    .A2(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5545_ (.A1(_1727_),
    .A2(_1729_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5546_ (.A1(\dspArea_regP[21] ),
    .A2(_1634_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5547_ (.A1(_1633_),
    .A2(_1635_),
    .B(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5548_ (.A1(_1726_),
    .A2(_1730_),
    .A3(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5549_ (.I(_1632_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5550_ (.A1(_1636_),
    .A2(_1638_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5551_ (.A1(_1636_),
    .A2(_1638_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5552_ (.A1(_1734_),
    .A2(_1735_),
    .B(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5553_ (.A1(_1733_),
    .A2(_1737_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5554_ (.A1(_1720_),
    .A2(_1738_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5555_ (.A1(_1642_),
    .A2(_1647_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5556_ (.A1(_1639_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5557_ (.A1(_1627_),
    .A2(_1644_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5558_ (.A1(_1741_),
    .A2(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5559_ (.A1(_1706_),
    .A2(_1739_),
    .A3(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5560_ (.A1(_1648_),
    .A2(_1649_),
    .A3(_1645_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5561_ (.A1(_1648_),
    .A2(_1649_),
    .B(_1645_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5562_ (.A1(_1613_),
    .A2(_1745_),
    .B(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5563_ (.A1(_1744_),
    .A2(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5564_ (.A1(_1682_),
    .A2(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5565_ (.A1(_1505_),
    .A2(_1541_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5566_ (.A1(_1652_),
    .A2(_1750_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5567_ (.A1(_1651_),
    .A2(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5568_ (.A1(_1589_),
    .A2(_1654_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5569_ (.A1(_1752_),
    .A2(_1753_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5570_ (.A1(_1667_),
    .A2(_1749_),
    .A3(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5571_ (.A1(_1655_),
    .A2(_1658_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5572_ (.A1(_1655_),
    .A2(_1658_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5573_ (.A1(_1574_),
    .A2(_1756_),
    .B(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5574_ (.A1(_1755_),
    .A2(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5575_ (.A1(_1574_),
    .A2(_1756_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5576_ (.A1(_1574_),
    .A2(_1756_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5577_ (.A1(_1571_),
    .A2(_1760_),
    .A3(_1761_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5578_ (.A1(_1465_),
    .A2(_1569_),
    .B(_1570_),
    .C(_1659_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5579_ (.A1(_1550_),
    .A2(_1552_),
    .A3(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5580_ (.A1(_1762_),
    .A2(_1764_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5581_ (.I(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5582_ (.A1(_1553_),
    .A2(_1554_),
    .A3(_1660_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5583_ (.A1(_1558_),
    .A2(_1559_),
    .A3(_1563_),
    .B(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5584_ (.A1(_1766_),
    .A2(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5585_ (.A1(_1759_),
    .A2(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5586_ (.I0(\dspArea_regP[22] ),
    .I1(_1770_),
    .S(_0441_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5587_ (.A1(_0355_),
    .A2(_1771_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5588_ (.A1(\dspArea_regP[23] ),
    .A2(_0259_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5589_ (.I(_0791_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5590_ (.A1(_1752_),
    .A2(_1753_),
    .A3(_1749_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5591_ (.A1(_1752_),
    .A2(_1753_),
    .B(_1749_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5592_ (.A1(_1667_),
    .A2(_1774_),
    .B(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5593_ (.A1(_1672_),
    .A2(_1680_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5594_ (.I(_1669_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5595_ (.A1(_1778_),
    .A2(_1681_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5596_ (.A1(_1777_),
    .A2(_1779_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5597_ (.A1(_0242_),
    .A2(_3034_),
    .A3(_1678_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5598_ (.A1(_1677_),
    .A2(_1781_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5599_ (.I(_1782_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5600_ (.A1(_1616_),
    .A2(_1626_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5601_ (.A1(_1625_),
    .A2(_1784_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5602_ (.A1(_1785_),
    .A2(_1702_),
    .B(_1705_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5603_ (.A1(_0228_),
    .A2(_3050_),
    .A3(_1598_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5604_ (.A1(_0233_),
    .A2(_3042_),
    .A3(_1692_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5605_ (.A1(_0236_),
    .A2(_3042_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5606_ (.A1(_1787_),
    .A2(_1788_),
    .A3(_1789_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5607_ (.A1(_1787_),
    .A2(_1788_),
    .B(_1789_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5608_ (.A1(_1790_),
    .A2(_1791_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5609_ (.A1(_0240_),
    .A2(_3038_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5610_ (.A1(_1792_),
    .A2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5611_ (.A1(_1786_),
    .A2(_1794_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5612_ (.A1(_1783_),
    .A2(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5613_ (.I(_1701_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5614_ (.A1(_1698_),
    .A2(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5615_ (.A1(_1698_),
    .A2(_1701_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5616_ (.A1(_1693_),
    .A2(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5617_ (.A1(_1710_),
    .A2(_1711_),
    .A3(_1716_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5618_ (.A1(_1709_),
    .A2(_1801_),
    .B(_1718_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5619_ (.A1(_0231_),
    .A2(_3045_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5620_ (.A1(_0225_),
    .A2(_3048_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5621_ (.A1(_0221_),
    .A2(_3052_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5622_ (.A1(_1804_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5623_ (.A1(_1803_),
    .A2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5624_ (.A1(_0216_),
    .A2(_3057_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5625_ (.A1(_0209_),
    .A2(_3060_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5626_ (.A1(_0205_),
    .A2(_3064_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5627_ (.A1(_1809_),
    .A2(_1810_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5628_ (.A1(_1808_),
    .A2(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5629_ (.A1(_0212_),
    .A2(_3061_),
    .A3(_1603_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5630_ (.A1(_0218_),
    .A2(_3053_),
    .A3(_1697_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5631_ (.A1(_1813_),
    .A2(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5632_ (.A1(_1807_),
    .A2(_1812_),
    .A3(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5633_ (.A1(_1802_),
    .A2(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5634_ (.A1(_1798_),
    .A2(_1800_),
    .A3(_1817_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5635_ (.A1(_1798_),
    .A2(_1800_),
    .B(_1817_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5636_ (.A1(_1818_),
    .A2(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5637_ (.A1(_0198_),
    .A2(_3076_),
    .A3(_1621_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5638_ (.A1(_0203_),
    .A2(_3066_),
    .A3(_1715_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5639_ (.A1(_1821_),
    .A2(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5640_ (.A1(_0184_),
    .A2(_3090_),
    .A3(_1630_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5641_ (.A1(_0190_),
    .A2(_3081_),
    .A3(_1724_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5642_ (.A1(_0201_),
    .A2(_3069_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5643_ (.A1(_0196_),
    .A2(_3075_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5644_ (.A1(_0193_),
    .A2(_3080_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5645_ (.A1(_1827_),
    .A2(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5646_ (.A1(_1826_),
    .A2(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5647_ (.A1(_1824_),
    .A2(_1825_),
    .A3(_1830_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5648_ (.A1(_1824_),
    .A2(_1825_),
    .B(_1830_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5649_ (.A1(_1831_),
    .A2(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5650_ (.A1(_1823_),
    .A2(_1833_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5651_ (.A1(_0188_),
    .A2(_3085_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5652_ (.A1(_0181_),
    .A2(_3089_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5653_ (.A1(_0176_),
    .A2(\dspArea_regA[21] ),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5654_ (.A1(_1836_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5655_ (.A1(_1835_),
    .A2(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5656_ (.I(_1839_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5657_ (.A1(_0172_),
    .A2(_3097_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5658_ (.A1(_0529_),
    .A2(_3101_),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5659_ (.A1(\dspArea_regP[23] ),
    .A2(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5660_ (.A1(_1841_),
    .A2(_1843_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5661_ (.A1(\dspArea_regP[22] ),
    .A2(_1728_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5662_ (.A1(_1727_),
    .A2(_1729_),
    .B(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5663_ (.A1(_1844_),
    .A2(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5664_ (.A1(_1840_),
    .A2(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5665_ (.A1(_1730_),
    .A2(_1732_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5666_ (.A1(_1730_),
    .A2(_1732_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5667_ (.A1(_1726_),
    .A2(_1849_),
    .B(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5668_ (.A1(_1848_),
    .A2(_1851_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5669_ (.A1(_1834_),
    .A2(_1852_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5670_ (.A1(_1733_),
    .A2(_1737_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5671_ (.A1(_1720_),
    .A2(_1738_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5672_ (.A1(_1854_),
    .A2(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5673_ (.A1(_1820_),
    .A2(_1853_),
    .A3(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5674_ (.A1(_1741_),
    .A2(_1742_),
    .A3(_1739_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5675_ (.A1(_1741_),
    .A2(_1742_),
    .B(_1739_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5676_ (.A1(_1706_),
    .A2(_1858_),
    .B(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5677_ (.A1(_1796_),
    .A2(_1857_),
    .A3(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5678_ (.A1(_1744_),
    .A2(_1747_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5679_ (.A1(_1682_),
    .A2(_1748_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5680_ (.A1(_1862_),
    .A2(_1863_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5681_ (.A1(_1780_),
    .A2(_1861_),
    .A3(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5682_ (.A1(_1776_),
    .A2(_1865_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5683_ (.A1(_1755_),
    .A2(_1758_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5684_ (.A1(_1755_),
    .A2(_1758_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5685_ (.A1(_1766_),
    .A2(_1768_),
    .B(_1868_),
    .C(_1867_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5686_ (.A1(_1867_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5687_ (.A1(_1866_),
    .A2(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5688_ (.A1(_1866_),
    .A2(_1870_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5689_ (.A1(_1773_),
    .A2(_1871_),
    .A3(_1872_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5690_ (.A1(_3173_),
    .A2(_1772_),
    .A3(_1873_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5691_ (.A1(_1786_),
    .A2(_1794_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5692_ (.A1(_1783_),
    .A2(_1795_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5693_ (.A1(_1874_),
    .A2(_1875_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5694_ (.A1(_0242_),
    .A2(_3038_),
    .A3(_1792_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5695_ (.A1(_1791_),
    .A2(_1877_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5696_ (.I(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5697_ (.A1(_1709_),
    .A2(_1719_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5698_ (.A1(_1718_),
    .A2(_1880_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5699_ (.A1(_1881_),
    .A2(_1816_),
    .B(_1819_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5700_ (.A1(_0228_),
    .A2(_3054_),
    .A3(_1691_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5701_ (.A1(_0233_),
    .A2(_3046_),
    .A3(_1806_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5702_ (.A1(_0236_),
    .A2(_3046_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5703_ (.A1(_1883_),
    .A2(_1884_),
    .A3(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5704_ (.A1(_1883_),
    .A2(_1884_),
    .B(_1885_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5705_ (.A1(_1886_),
    .A2(_1887_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5706_ (.A1(_0240_),
    .A2(_3042_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5707_ (.A1(_1888_),
    .A2(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5708_ (.A1(_1882_),
    .A2(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5709_ (.A1(_1879_),
    .A2(_1891_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5710_ (.I(_1815_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5711_ (.A1(_1812_),
    .A2(_1893_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5712_ (.A1(_1812_),
    .A2(_1815_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5713_ (.A1(_1807_),
    .A2(_1895_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5714_ (.A1(_1824_),
    .A2(_1825_),
    .A3(_1830_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5715_ (.A1(_1823_),
    .A2(_1897_),
    .B(_1832_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5716_ (.A1(_0232_),
    .A2(_3049_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5717_ (.A1(_0226_),
    .A2(_3052_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5718_ (.A1(_0222_),
    .A2(_3056_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5719_ (.A1(_1900_),
    .A2(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5720_ (.A1(_1899_),
    .A2(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5721_ (.A1(_0217_),
    .A2(_3061_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5722_ (.A1(_0210_),
    .A2(_3064_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5723_ (.A1(_0206_),
    .A2(_3068_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5724_ (.A1(_1905_),
    .A2(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5725_ (.A1(_1904_),
    .A2(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5726_ (.A1(_0213_),
    .A2(_3065_),
    .A3(_1696_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5727_ (.A1(_0219_),
    .A2(_3057_),
    .A3(_1811_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5728_ (.A1(_1909_),
    .A2(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5729_ (.A1(_1903_),
    .A2(_1908_),
    .A3(_1911_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5730_ (.A1(_1898_),
    .A2(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5731_ (.A1(_1894_),
    .A2(_1896_),
    .A3(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5732_ (.A1(_1894_),
    .A2(_1896_),
    .B(_1913_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5733_ (.A1(_1914_),
    .A2(_1915_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5734_ (.A1(_0197_),
    .A2(_3081_),
    .A3(_1714_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5735_ (.A1(_0202_),
    .A2(_3070_),
    .A3(_1829_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5736_ (.A1(_1917_),
    .A2(_1918_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5737_ (.A1(_0183_),
    .A2(_3093_),
    .A3(_1723_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5738_ (.A1(_0189_),
    .A2(_3086_),
    .A3(_1838_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5739_ (.A1(_0404_),
    .A2(_3075_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5740_ (.A1(_0364_),
    .A2(_3079_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5741_ (.A1(_0406_),
    .A2(_3084_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5742_ (.A1(_1923_),
    .A2(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5743_ (.A1(_1922_),
    .A2(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5744_ (.A1(_1920_),
    .A2(_1921_),
    .A3(_1926_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5745_ (.A1(_1920_),
    .A2(_1921_),
    .B(_1926_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5746_ (.A1(_1927_),
    .A2(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5747_ (.A1(_1919_),
    .A2(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5748_ (.A1(_0187_),
    .A2(_3089_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5749_ (.A1(_0180_),
    .A2(\dspArea_regA[21] ),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5750_ (.A1(_0176_),
    .A2(\dspArea_regA[22] ),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5751_ (.A1(_1932_),
    .A2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5752_ (.A1(_1931_),
    .A2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5753_ (.A1(_0173_),
    .A2(_3101_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5754_ (.A1(_0167_),
    .A2(\dspArea_regA[24] ),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5755_ (.A1(\dspArea_regP[24] ),
    .A2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5756_ (.A1(_1936_),
    .A2(_1938_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5757_ (.A1(\dspArea_regP[23] ),
    .A2(_1842_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5758_ (.A1(_1841_),
    .A2(_1843_),
    .B(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5759_ (.A1(_1935_),
    .A2(_1939_),
    .A3(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5760_ (.A1(_1844_),
    .A2(_1846_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5761_ (.A1(_1844_),
    .A2(_1846_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5762_ (.A1(_1840_),
    .A2(_1943_),
    .B(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5763_ (.A1(_1942_),
    .A2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5764_ (.A1(_1930_),
    .A2(_1946_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5765_ (.A1(_1848_),
    .A2(_1851_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5766_ (.A1(_1834_),
    .A2(_1852_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5767_ (.A1(_1948_),
    .A2(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5768_ (.A1(_1916_),
    .A2(_1947_),
    .A3(_1950_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5769_ (.A1(_1854_),
    .A2(_1855_),
    .A3(_1853_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5770_ (.A1(_1854_),
    .A2(_1855_),
    .B(_1853_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5771_ (.A1(_1820_),
    .A2(_1952_),
    .B(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5772_ (.A1(_1892_),
    .A2(_1951_),
    .A3(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5773_ (.A1(_1857_),
    .A2(_1860_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5774_ (.A1(_1857_),
    .A2(_1860_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5775_ (.A1(_1796_),
    .A2(_1956_),
    .B(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5776_ (.A1(_1955_),
    .A2(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5777_ (.A1(_1876_),
    .A2(_1959_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5778_ (.A1(_1862_),
    .A2(_1863_),
    .A3(_1861_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5779_ (.A1(_1862_),
    .A2(_1863_),
    .B(_1861_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5780_ (.A1(_1780_),
    .A2(_1961_),
    .B(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5781_ (.A1(_1960_),
    .A2(_1963_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5782_ (.I(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5783_ (.A1(_1759_),
    .A2(_1866_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5784_ (.A1(_1558_),
    .A2(_1559_),
    .B(_1767_),
    .C(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5785_ (.A1(_1776_),
    .A2(_1865_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5786_ (.A1(_1867_),
    .A2(_1968_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5787_ (.A1(_1776_),
    .A2(_1865_),
    .B1(_1966_),
    .B2(_1765_),
    .C(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5788_ (.A1(_1967_),
    .A2(_1970_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5789_ (.A1(_1159_),
    .A2(_1252_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _5790_ (.A1(_1972_),
    .A2(_1561_),
    .A3(_1767_),
    .A4(_1966_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5791_ (.A1(_1257_),
    .A2(_1258_),
    .B(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5792_ (.A1(_1971_),
    .A2(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5793_ (.A1(_1965_),
    .A2(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5794_ (.I0(\dspArea_regP[24] ),
    .I1(_1976_),
    .S(_0441_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5795_ (.A1(_0355_),
    .A2(_1977_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5796_ (.I(\dspArea_regP[25] ),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5797_ (.A1(_1955_),
    .A2(_1958_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5798_ (.A1(_1876_),
    .A2(_1959_),
    .B(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5799_ (.A1(_1882_),
    .A2(_1890_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5800_ (.A1(_1879_),
    .A2(_1891_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5801_ (.A1(_1981_),
    .A2(_1982_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5802_ (.A1(_0244_),
    .A2(_3042_),
    .A3(_1888_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5803_ (.A1(_1887_),
    .A2(_1984_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5804_ (.A1(_1823_),
    .A2(_1833_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5805_ (.A1(_1832_),
    .A2(_1986_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5806_ (.A1(_1987_),
    .A2(_1912_),
    .B(_1915_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5807_ (.A1(_0229_),
    .A2(_3058_),
    .A3(_1805_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5808_ (.A1(_0234_),
    .A2(_3050_),
    .A3(_1902_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5809_ (.A1(_0237_),
    .A2(_3050_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5810_ (.A1(_1989_),
    .A2(_1990_),
    .A3(_1991_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5811_ (.A1(_1989_),
    .A2(_1990_),
    .B(_1991_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5812_ (.A1(_1992_),
    .A2(_1993_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5813_ (.A1(_0242_),
    .A2(_3046_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5814_ (.A1(_1994_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5815_ (.A1(_1988_),
    .A2(_1996_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5816_ (.A1(_1985_),
    .A2(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5817_ (.I(_1911_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5818_ (.A1(_1908_),
    .A2(_1999_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5819_ (.A1(_1908_),
    .A2(_1911_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5820_ (.A1(_1903_),
    .A2(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5821_ (.A1(_1920_),
    .A2(_1921_),
    .A3(_1926_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5822_ (.A1(_1919_),
    .A2(_2003_),
    .B(_1928_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5823_ (.A1(_0231_),
    .A2(_3053_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5824_ (.A1(_0226_),
    .A2(_3056_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5825_ (.A1(_0221_),
    .A2(_3060_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5826_ (.A1(_2006_),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5827_ (.A1(_2005_),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5828_ (.A1(_0216_),
    .A2(_3065_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5829_ (.A1(_0210_),
    .A2(_3068_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5830_ (.A1(_0206_),
    .A2(_3074_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5831_ (.A1(_2011_),
    .A2(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5832_ (.A1(_2010_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5833_ (.A1(_0212_),
    .A2(_3069_),
    .A3(_1810_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5834_ (.A1(_0634_),
    .A2(_3061_),
    .A3(_1907_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5835_ (.A1(_2015_),
    .A2(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5836_ (.A1(_2009_),
    .A2(_2014_),
    .A3(_2017_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5837_ (.A1(_2004_),
    .A2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5838_ (.A1(_2000_),
    .A2(_2002_),
    .A3(_2019_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5839_ (.A1(_2000_),
    .A2(_2002_),
    .B(_2019_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5840_ (.A1(_2020_),
    .A2(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5841_ (.A1(_0197_),
    .A2(_3085_),
    .A3(_1828_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5842_ (.A1(_0202_),
    .A2(_3076_),
    .A3(_1925_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5843_ (.A1(_2023_),
    .A2(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5844_ (.A1(_0183_),
    .A2(_3097_),
    .A3(_1837_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5845_ (.A1(_0188_),
    .A2(_3090_),
    .A3(_1934_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5846_ (.A1(_0404_),
    .A2(_3080_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5847_ (.A1(_0195_),
    .A2(_3084_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5848_ (.A1(_0192_),
    .A2(\dspArea_regA[20] ),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5849_ (.A1(_2029_),
    .A2(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5850_ (.A1(_2028_),
    .A2(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5851_ (.A1(_2026_),
    .A2(_2027_),
    .A3(_2032_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5852_ (.A1(_2026_),
    .A2(_2027_),
    .B(_2032_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5853_ (.A1(_2033_),
    .A2(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5854_ (.A1(_2025_),
    .A2(_2035_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5855_ (.A1(_0188_),
    .A2(_3093_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5856_ (.A1(_0181_),
    .A2(_3097_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5857_ (.A1(_0177_),
    .A2(_3101_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5858_ (.A1(_2038_),
    .A2(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5859_ (.A1(_2037_),
    .A2(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5860_ (.A1(_0172_),
    .A2(\dspArea_regA[24] ),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5861_ (.A1(_1978_),
    .A2(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5862_ (.A1(\dspArea_regP[24] ),
    .A2(_0168_),
    .A3(\dspArea_regA[24] ),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5863_ (.I(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5864_ (.A1(_1936_),
    .A2(_1938_),
    .B(_2045_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5865_ (.A1(_2043_),
    .A2(_2046_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5866_ (.A1(_2041_),
    .A2(_2047_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5867_ (.I(_1935_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5868_ (.A1(_1939_),
    .A2(_1941_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5869_ (.A1(_1939_),
    .A2(_1941_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5870_ (.A1(_2049_),
    .A2(_2050_),
    .B(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5871_ (.A1(_2048_),
    .A2(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5872_ (.A1(_2036_),
    .A2(_2053_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5873_ (.A1(_1839_),
    .A2(_1847_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5874_ (.A1(_1944_),
    .A2(_2055_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5875_ (.A1(_1942_),
    .A2(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5876_ (.A1(_1930_),
    .A2(_1946_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5877_ (.A1(_2057_),
    .A2(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5878_ (.A1(_2022_),
    .A2(_2054_),
    .A3(_2059_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5879_ (.A1(_1948_),
    .A2(_1949_),
    .A3(_1947_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5880_ (.A1(_1948_),
    .A2(_1949_),
    .B(_1947_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5881_ (.A1(_1916_),
    .A2(_2061_),
    .B(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5882_ (.A1(_2060_),
    .A2(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5883_ (.A1(_1998_),
    .A2(_2064_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5884_ (.A1(_1951_),
    .A2(_1954_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5885_ (.A1(_1951_),
    .A2(_1954_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5886_ (.A1(_1892_),
    .A2(_2066_),
    .B(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5887_ (.A1(_1983_),
    .A2(_2065_),
    .A3(_2068_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5888_ (.A1(_1980_),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5889_ (.A1(_1960_),
    .A2(_1963_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5890_ (.A1(_1964_),
    .A2(_1975_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5891_ (.A1(_2071_),
    .A2(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5892_ (.A1(_2070_),
    .A2(_2073_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5893_ (.A1(_1773_),
    .A2(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5894_ (.A1(_1978_),
    .A2(_0297_),
    .B(_2075_),
    .C(_1461_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5895_ (.I(\dspArea_regP[26] ),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5896_ (.A1(_1988_),
    .A2(_1996_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5897_ (.I(_1985_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5898_ (.A1(_2078_),
    .A2(_1997_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5899_ (.A1(_2077_),
    .A2(_2079_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5900_ (.A1(_0243_),
    .A2(_3046_),
    .A3(_1994_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5901_ (.A1(_1993_),
    .A2(_2081_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5902_ (.I(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5903_ (.A1(_1919_),
    .A2(_1929_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5904_ (.A1(_1928_),
    .A2(_2084_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5905_ (.A1(_2085_),
    .A2(_2018_),
    .B(_2021_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5906_ (.A1(_0228_),
    .A2(_3062_),
    .A3(_1901_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5907_ (.A1(_0233_),
    .A2(_3054_),
    .A3(_2008_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5908_ (.A1(_0236_),
    .A2(_3054_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5909_ (.A1(_2087_),
    .A2(_2088_),
    .A3(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5910_ (.A1(_2087_),
    .A2(_2088_),
    .B(_2089_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5911_ (.A1(_2090_),
    .A2(_2091_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5912_ (.A1(_0240_),
    .A2(_3050_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5913_ (.A1(_2092_),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5914_ (.A1(_2086_),
    .A2(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5915_ (.A1(_2083_),
    .A2(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5916_ (.I(_2017_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5917_ (.A1(_2014_),
    .A2(_2097_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5918_ (.A1(_2014_),
    .A2(_2017_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5919_ (.A1(_2009_),
    .A2(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5920_ (.A1(_2026_),
    .A2(_2027_),
    .A3(_2032_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5921_ (.A1(_2025_),
    .A2(_2101_),
    .B(_2034_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5922_ (.A1(\dspArea_regB[13] ),
    .A2(_3057_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5923_ (.A1(_0225_),
    .A2(_3060_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5924_ (.A1(\dspArea_regB[11] ),
    .A2(_3064_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5925_ (.A1(_2104_),
    .A2(_2105_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5926_ (.A1(_2103_),
    .A2(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5927_ (.A1(_0216_),
    .A2(_3069_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5928_ (.A1(_0209_),
    .A2(_3074_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5929_ (.A1(_0205_),
    .A2(_3079_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5930_ (.A1(_2109_),
    .A2(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5931_ (.A1(_2108_),
    .A2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5932_ (.A1(_0211_),
    .A2(_3075_),
    .A3(_1906_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5933_ (.A1(_0217_),
    .A2(_3065_),
    .A3(_2013_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5934_ (.A1(_2113_),
    .A2(_2114_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5935_ (.A1(_2107_),
    .A2(_2112_),
    .A3(_2115_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5936_ (.A1(_2102_),
    .A2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5937_ (.A1(_2098_),
    .A2(_2100_),
    .A3(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5938_ (.A1(_2098_),
    .A2(_2100_),
    .B(_2117_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5939_ (.A1(_2118_),
    .A2(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5940_ (.A1(_0198_),
    .A2(_3090_),
    .A3(_1924_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5941_ (.A1(_0202_),
    .A2(_3081_),
    .A3(_2031_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5942_ (.A1(_2121_),
    .A2(_2122_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5943_ (.A1(_0181_),
    .A2(_3101_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5944_ (.A1(_1933_),
    .A2(_2124_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5945_ (.A1(_0188_),
    .A2(_3093_),
    .A3(_2040_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5946_ (.A1(_0404_),
    .A2(_3085_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5947_ (.A1(_0195_),
    .A2(\dspArea_regA[20] ),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5948_ (.A1(_0192_),
    .A2(\dspArea_regA[21] ),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5949_ (.A1(_2128_),
    .A2(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5950_ (.A1(_2127_),
    .A2(_2130_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5951_ (.A1(_2125_),
    .A2(_2126_),
    .A3(_2131_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5952_ (.A1(_2125_),
    .A2(_2126_),
    .B(_2131_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5953_ (.A1(_2132_),
    .A2(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5954_ (.A1(_2123_),
    .A2(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5955_ (.A1(\dspArea_regP[25] ),
    .A2(_0173_),
    .A3(_3105_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5956_ (.A1(\dspArea_regP[26] ),
    .A2(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5957_ (.A1(_0186_),
    .A2(_3097_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5958_ (.A1(_0177_),
    .A2(_3105_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5959_ (.A1(_2124_),
    .A2(_2138_),
    .A3(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5960_ (.A1(_2137_),
    .A2(_2140_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5961_ (.A1(_2043_),
    .A2(_2046_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5962_ (.A1(_2041_),
    .A2(_2047_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5963_ (.A1(_2142_),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5964_ (.A1(_2135_),
    .A2(_2141_),
    .A3(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5965_ (.A1(_2048_),
    .A2(_2052_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5966_ (.A1(_2036_),
    .A2(_2053_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5967_ (.A1(_2146_),
    .A2(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5968_ (.A1(_2120_),
    .A2(_2145_),
    .A3(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5969_ (.A1(_2057_),
    .A2(_2058_),
    .A3(_2054_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5970_ (.A1(_2057_),
    .A2(_2058_),
    .B(_2054_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5971_ (.A1(_2022_),
    .A2(_2150_),
    .B(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5972_ (.A1(_2096_),
    .A2(_2149_),
    .A3(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5973_ (.A1(_2060_),
    .A2(_2063_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5974_ (.A1(_1998_),
    .A2(_2064_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5975_ (.A1(_2154_),
    .A2(_2155_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _5976_ (.A1(_2080_),
    .A2(_2153_),
    .A3(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _5977_ (.A1(_2065_),
    .A2(_2068_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5978_ (.A1(_2065_),
    .A2(_2068_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _5979_ (.A1(_1983_),
    .A2(_2158_),
    .B(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5980_ (.A1(_2157_),
    .A2(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _5981_ (.A1(_1983_),
    .A2(_2158_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5982_ (.A1(_1983_),
    .A2(_2158_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5983_ (.A1(_1980_),
    .A2(_2162_),
    .A3(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5984_ (.A1(_1876_),
    .A2(_1959_),
    .B(_2069_),
    .C(_1979_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5985_ (.A1(_1960_),
    .A2(_1963_),
    .A3(_2165_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5986_ (.A1(_2164_),
    .A2(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5987_ (.I(_2070_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5988_ (.A1(_1971_),
    .A2(_1974_),
    .B(_2168_),
    .C(_1965_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _5989_ (.A1(_2161_),
    .A2(_2167_),
    .A3(_2169_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5990_ (.A1(_2167_),
    .A2(_2169_),
    .B(_2161_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5991_ (.A1(_2170_),
    .A2(_2171_),
    .B(_0248_),
    .C(_0790_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5992_ (.A1(_2076_),
    .A2(_0297_),
    .B(_2172_),
    .C(_1461_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5993_ (.I(\dspArea_regP[27] ),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5994_ (.A1(_2154_),
    .A2(_2155_),
    .A3(_2153_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5995_ (.A1(_2154_),
    .A2(_2155_),
    .B(_2153_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5996_ (.A1(_2080_),
    .A2(_2174_),
    .B(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5997_ (.A1(_2086_),
    .A2(_2094_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5998_ (.A1(_2083_),
    .A2(_2095_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5999_ (.A1(_2177_),
    .A2(_2178_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6000_ (.A1(_0242_),
    .A2(_3050_),
    .A3(_2092_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6001_ (.A1(_2091_),
    .A2(_2180_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6002_ (.I(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6003_ (.A1(_2025_),
    .A2(_2035_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6004_ (.A1(_2034_),
    .A2(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6005_ (.A1(_2184_),
    .A2(_2116_),
    .B(_2119_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6006_ (.A1(_0225_),
    .A2(_3064_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6007_ (.A1(_2007_),
    .A2(_2186_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6008_ (.A1(_0233_),
    .A2(_3058_),
    .A3(_2106_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6009_ (.A1(\dspArea_regB[14] ),
    .A2(_3058_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6010_ (.A1(_2187_),
    .A2(_2188_),
    .A3(_2189_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6011_ (.A1(_2187_),
    .A2(_2188_),
    .B(_2189_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6012_ (.A1(_2190_),
    .A2(_2191_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6013_ (.A1(_0240_),
    .A2(_3054_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6014_ (.A1(_2192_),
    .A2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6015_ (.A1(_2185_),
    .A2(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6016_ (.A1(_2182_),
    .A2(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6017_ (.I(_2115_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6018_ (.A1(_2112_),
    .A2(_2197_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6019_ (.A1(_2112_),
    .A2(_2115_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6020_ (.A1(_2107_),
    .A2(_2199_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6021_ (.A1(_2125_),
    .A2(_2126_),
    .A3(_2131_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6022_ (.A1(_2123_),
    .A2(_2201_),
    .B(_2133_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6023_ (.A1(_0231_),
    .A2(_3061_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6024_ (.A1(_0221_),
    .A2(_3068_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6025_ (.A1(_2186_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6026_ (.A1(_2203_),
    .A2(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6027_ (.A1(_0216_),
    .A2(_3075_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6028_ (.A1(_0210_),
    .A2(_3079_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6029_ (.A1(_0206_),
    .A2(_3084_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6030_ (.A1(_2208_),
    .A2(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6031_ (.A1(_2207_),
    .A2(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6032_ (.A1(_0212_),
    .A2(_3080_),
    .A3(_2012_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6033_ (.A1(_0634_),
    .A2(_3069_),
    .A3(_2111_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6034_ (.A1(_2212_),
    .A2(_2213_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6035_ (.A1(_2206_),
    .A2(_2211_),
    .A3(_2214_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6036_ (.A1(_2202_),
    .A2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6037_ (.A1(_2198_),
    .A2(_2200_),
    .A3(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6038_ (.A1(_2198_),
    .A2(_2200_),
    .B(_2216_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6039_ (.A1(_2217_),
    .A2(_2218_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6040_ (.A1(_0182_),
    .A2(_3105_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6041_ (.A1(_0188_),
    .A2(_3101_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6042_ (.A1(_2220_),
    .A2(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6043_ (.A1(_0187_),
    .A2(_3105_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6044_ (.A1(_2124_),
    .A2(_2223_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6045_ (.A1(_2222_),
    .A2(_2224_),
    .B(_2173_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6046_ (.A1(_2173_),
    .A2(_2222_),
    .A3(_2224_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6047_ (.A1(_2225_),
    .A2(_2226_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6048_ (.A1(\dspArea_regP[26] ),
    .A2(_2136_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6049_ (.A1(_2137_),
    .A2(_2140_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6050_ (.A1(_2228_),
    .A2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6051_ (.A1(_2227_),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6052_ (.A1(_0195_),
    .A2(\dspArea_regA[21] ),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6053_ (.A1(_2030_),
    .A2(_2232_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6054_ (.A1(_0202_),
    .A2(_3086_),
    .A3(_2130_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6055_ (.A1(_2233_),
    .A2(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6056_ (.I(_2138_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6057_ (.A1(_2124_),
    .A2(_2139_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6058_ (.A1(_0178_),
    .A2(_3105_),
    .A3(_2124_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6059_ (.A1(_2236_),
    .A2(_2237_),
    .B(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6060_ (.A1(_0200_),
    .A2(_3089_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6061_ (.A1(_0193_),
    .A2(_3097_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6062_ (.A1(_2232_),
    .A2(_2240_),
    .A3(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6063_ (.A1(_2239_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6064_ (.A1(_2235_),
    .A2(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6065_ (.A1(_2231_),
    .A2(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6066_ (.A1(_2142_),
    .A2(_2143_),
    .A3(_2141_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6067_ (.A1(_2142_),
    .A2(_2143_),
    .B(_2141_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6068_ (.A1(_2135_),
    .A2(_2246_),
    .B(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6069_ (.A1(_2245_),
    .A2(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6070_ (.A1(_2219_),
    .A2(_2249_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6071_ (.A1(_2146_),
    .A2(_2147_),
    .A3(_2145_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6072_ (.A1(_2146_),
    .A2(_2147_),
    .B(_2145_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6073_ (.A1(_2120_),
    .A2(_2251_),
    .B(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6074_ (.A1(_2196_),
    .A2(_2250_),
    .A3(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6075_ (.A1(_2149_),
    .A2(_2152_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6076_ (.A1(_2149_),
    .A2(_2152_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6077_ (.A1(_2096_),
    .A2(_2255_),
    .B(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6078_ (.A1(_2254_),
    .A2(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6079_ (.A1(_2179_),
    .A2(_2258_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6080_ (.A1(_2176_),
    .A2(_2259_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6081_ (.A1(_2157_),
    .A2(_2160_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6082_ (.A1(_2261_),
    .A2(_2171_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6083_ (.A1(_2260_),
    .A2(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6084_ (.A1(_2260_),
    .A2(_2262_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6085_ (.A1(_0296_),
    .A2(_2263_),
    .A3(_2264_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6086_ (.A1(_2173_),
    .A2(_0297_),
    .B(_2265_),
    .C(_1461_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6087_ (.A1(_2185_),
    .A2(_2194_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6088_ (.A1(_2182_),
    .A2(_2195_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6089_ (.A1(_2266_),
    .A2(_2267_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6090_ (.A1(_0243_),
    .A2(_3054_),
    .A3(_2192_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6091_ (.A1(_2191_),
    .A2(_2269_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6092_ (.I(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6093_ (.A1(_2123_),
    .A2(_2134_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6094_ (.A1(_2133_),
    .A2(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6095_ (.A1(_2273_),
    .A2(_2215_),
    .B(_2218_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6096_ (.A1(_0223_),
    .A2(_3070_),
    .A3(_2186_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6097_ (.A1(_0233_),
    .A2(_3062_),
    .A3(_2205_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6098_ (.A1(_0236_),
    .A2(_3062_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6099_ (.A1(_2275_),
    .A2(_2276_),
    .A3(_2277_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6100_ (.A1(_2275_),
    .A2(_2276_),
    .B(_2277_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6101_ (.A1(_2278_),
    .A2(_2279_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6102_ (.A1(_0240_),
    .A2(_3058_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6103_ (.A1(_2280_),
    .A2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6104_ (.A1(_2274_),
    .A2(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6105_ (.A1(_2271_),
    .A2(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6106_ (.A1(\dspArea_regP[28] ),
    .A2(_2223_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6107_ (.A1(_2232_),
    .A2(_2241_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6108_ (.A1(_0196_),
    .A2(_3097_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6109_ (.A1(_2129_),
    .A2(_2287_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6110_ (.A1(_2240_),
    .A2(_2286_),
    .B(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6111_ (.A1(_0200_),
    .A2(_3093_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6112_ (.A1(_0193_),
    .A2(_3101_),
    .Z(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6113_ (.A1(_2287_),
    .A2(_2290_),
    .A3(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6114_ (.A1(_2224_),
    .A2(_2292_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6115_ (.A1(_2289_),
    .A2(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6116_ (.A1(_2226_),
    .A2(_2285_),
    .A3(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6117_ (.A1(_2228_),
    .A2(_2229_),
    .B(_2227_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6118_ (.I(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6119_ (.A1(_2231_),
    .A2(_2244_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6120_ (.A1(_2297_),
    .A2(_2298_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6121_ (.A1(_2212_),
    .A2(_2213_),
    .B(_2211_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6122_ (.A1(_2212_),
    .A2(_2213_),
    .A3(_2211_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6123_ (.A1(_2206_),
    .A2(_2301_),
    .A3(_2300_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6124_ (.A1(_2300_),
    .A2(_2302_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6125_ (.A1(_2239_),
    .A2(_2242_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6126_ (.I(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6127_ (.A1(_2235_),
    .A2(_2243_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6128_ (.A1(_2305_),
    .A2(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6129_ (.A1(_0232_),
    .A2(_3066_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6130_ (.A1(_0227_),
    .A2(_3069_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6131_ (.A1(_0222_),
    .A2(_3075_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6132_ (.A1(_2309_),
    .A2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6133_ (.A1(_2308_),
    .A2(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6134_ (.A1(_0212_),
    .A2(_3085_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6135_ (.A1(_0634_),
    .A2(_3080_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6136_ (.A1(_0207_),
    .A2(_3089_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6137_ (.A1(_2313_),
    .A2(_2314_),
    .A3(_2315_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6138_ (.A1(_0213_),
    .A2(_3086_),
    .A3(_2110_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6139_ (.A1(_0219_),
    .A2(_3076_),
    .A3(_2210_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6140_ (.A1(_2317_),
    .A2(_2318_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6141_ (.A1(_2312_),
    .A2(_2316_),
    .A3(_2319_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6142_ (.A1(_2303_),
    .A2(_2307_),
    .A3(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6143_ (.A1(_2295_),
    .A2(_2299_),
    .A3(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6144_ (.I(_2245_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6145_ (.A1(_2323_),
    .A2(_2248_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6146_ (.A1(_2219_),
    .A2(_2249_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6147_ (.A1(_2324_),
    .A2(_2325_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6148_ (.A1(_2284_),
    .A2(_2322_),
    .A3(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6149_ (.A1(_2250_),
    .A2(_2253_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6150_ (.A1(_2250_),
    .A2(_2253_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6151_ (.A1(_2196_),
    .A2(_2328_),
    .B(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6152_ (.A1(_2327_),
    .A2(_2330_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6153_ (.A1(_2254_),
    .A2(_2257_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6154_ (.A1(_2179_),
    .A2(_2258_),
    .B(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6155_ (.A1(_2268_),
    .A2(_2331_),
    .A3(_2333_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6156_ (.A1(_2176_),
    .A2(_2259_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6157_ (.A1(_2157_),
    .A2(_2160_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6158_ (.A1(_2164_),
    .A2(_2166_),
    .B(_2335_),
    .C(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6159_ (.A1(_2176_),
    .A2(_2259_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6160_ (.A1(_2176_),
    .A2(_2259_),
    .B(_2157_),
    .C(_2160_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6161_ (.A1(_2338_),
    .A2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6162_ (.A1(_1964_),
    .A2(_2070_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6163_ (.A1(_2161_),
    .A2(_2260_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6164_ (.A1(_1971_),
    .A2(_1974_),
    .B(_2341_),
    .C(_2342_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6165_ (.A1(_2337_),
    .A2(_2340_),
    .A3(_2343_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6166_ (.A1(_2334_),
    .A2(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6167_ (.I0(\dspArea_regP[28] ),
    .I1(_2345_),
    .S(_0441_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6168_ (.A1(_3111_),
    .A2(_2346_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6169_ (.A1(_2327_),
    .A2(_2330_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6170_ (.A1(_2268_),
    .A2(_2331_),
    .B(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6171_ (.A1(_2274_),
    .A2(_2282_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6172_ (.A1(_2271_),
    .A2(_2283_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6173_ (.A1(_2349_),
    .A2(_2350_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6174_ (.A1(\dspArea_regP[28] ),
    .A2(_2223_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6175_ (.A1(\dspArea_regP[29] ),
    .A2(_2352_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6176_ (.A1(_0201_),
    .A2(_3097_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6177_ (.A1(_0196_),
    .A2(_3101_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6178_ (.A1(_0193_),
    .A2(\dspArea_regA[24] ),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6179_ (.A1(_2355_),
    .A2(_2356_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6180_ (.A1(_2354_),
    .A2(_2357_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6181_ (.A1(_2287_),
    .A2(_2291_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6182_ (.A1(_2241_),
    .A2(_2355_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6183_ (.A1(_2290_),
    .A2(_2359_),
    .B(_2360_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6184_ (.A1(_2358_),
    .A2(_2361_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6185_ (.A1(_2353_),
    .A2(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6186_ (.A1(_2226_),
    .A2(_2285_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6187_ (.A1(_2226_),
    .A2(_2285_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6188_ (.A1(_2364_),
    .A2(_2294_),
    .B(_2365_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6189_ (.A1(_2363_),
    .A2(_2366_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6190_ (.A1(_2317_),
    .A2(_2318_),
    .A3(_2316_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6191_ (.A1(_2317_),
    .A2(_2318_),
    .B(_2316_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6192_ (.A1(_2312_),
    .A2(_2368_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6193_ (.A1(_2224_),
    .A2(_2292_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6194_ (.A1(_2289_),
    .A2(_2293_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6195_ (.A1(_2371_),
    .A2(_2372_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6196_ (.A1(_0232_),
    .A2(_3070_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6197_ (.A1(_0227_),
    .A2(_3075_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6198_ (.A1(_0223_),
    .A2(_3080_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6199_ (.A1(_2375_),
    .A2(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6200_ (.A1(_2374_),
    .A2(_2377_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6201_ (.A1(_0218_),
    .A2(_3085_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6202_ (.A1(_0211_),
    .A2(_3089_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6203_ (.A1(_0207_),
    .A2(_3093_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6204_ (.A1(_2380_),
    .A2(_2381_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6205_ (.A1(_2379_),
    .A2(_2382_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6206_ (.A1(_2313_),
    .A2(_2315_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6207_ (.A1(_2209_),
    .A2(_2380_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6208_ (.A1(_2314_),
    .A2(_2384_),
    .B(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6209_ (.A1(_2383_),
    .A2(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6210_ (.A1(_2378_),
    .A2(_2387_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6211_ (.A1(_2370_),
    .A2(_2373_),
    .A3(_2388_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6212_ (.A1(_2367_),
    .A2(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6213_ (.I(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6214_ (.A1(_2297_),
    .A2(_2298_),
    .A3(_2295_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6215_ (.A1(_2297_),
    .A2(_2298_),
    .B(_2295_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6216_ (.A1(_2392_),
    .A2(_2321_),
    .B(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6217_ (.A1(_0244_),
    .A2(_3058_),
    .A3(_2280_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6218_ (.A1(_2279_),
    .A2(_2395_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6219_ (.A1(_2305_),
    .A2(_2306_),
    .A3(_2320_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6220_ (.A1(_2305_),
    .A2(_2306_),
    .B(_2320_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6221_ (.A1(_2303_),
    .A2(_2397_),
    .B(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6222_ (.A1(_2308_),
    .A2(_2311_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6223_ (.A1(_2204_),
    .A2(_2375_),
    .B(_2400_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6224_ (.A1(_0237_),
    .A2(_3066_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6225_ (.A1(_2401_),
    .A2(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6226_ (.A1(_0241_),
    .A2(_3062_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6227_ (.A1(_2403_),
    .A2(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6228_ (.A1(_2399_),
    .A2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6229_ (.A1(_2396_),
    .A2(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6230_ (.A1(_2391_),
    .A2(_2394_),
    .A3(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6231_ (.A1(_2324_),
    .A2(_2325_),
    .A3(_2322_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6232_ (.A1(_2324_),
    .A2(_2325_),
    .B(_2322_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6233_ (.A1(_2284_),
    .A2(_2409_),
    .B(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6234_ (.A1(_2351_),
    .A2(_2408_),
    .A3(_2411_),
    .Z(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6235_ (.A1(_2348_),
    .A2(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6236_ (.I(_2334_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6237_ (.A1(_2268_),
    .A2(_2331_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6238_ (.A1(_2268_),
    .A2(_2331_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6239_ (.A1(_2415_),
    .A2(_2416_),
    .A3(_2333_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6240_ (.A1(_2414_),
    .A2(_2344_),
    .B(_2417_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6241_ (.A1(_2413_),
    .A2(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6242_ (.A1(\dspArea_regP[29] ),
    .A2(_0874_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6243_ (.A1(_0792_),
    .A2(_2419_),
    .B(_2420_),
    .C(_1461_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6244_ (.A1(_0197_),
    .A2(_3105_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6245_ (.A1(_0202_),
    .A2(_3102_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6246_ (.A1(_2421_),
    .A2(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6247_ (.A1(_2421_),
    .A2(_2422_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6248_ (.A1(_2423_),
    .A2(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6249_ (.A1(_0193_),
    .A2(_3105_),
    .A3(_2355_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6250_ (.A1(_2354_),
    .A2(_2357_),
    .B(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6251_ (.A1(_2425_),
    .A2(_2427_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6252_ (.A1(\dspArea_regP[30] ),
    .A2(_2428_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6253_ (.A1(\dspArea_regP[29] ),
    .A2(_2352_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6254_ (.A1(_2353_),
    .A2(_2362_),
    .B(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6255_ (.A1(_2429_),
    .A2(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6256_ (.I(_2378_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6257_ (.A1(_2383_),
    .A2(_2386_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6258_ (.A1(_2433_),
    .A2(_2387_),
    .B(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6259_ (.A1(_2358_),
    .A2(_2361_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6260_ (.A1(_0232_),
    .A2(_3075_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6261_ (.A1(_0226_),
    .A2(_3080_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6262_ (.A1(_0222_),
    .A2(_3085_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6263_ (.A1(_2438_),
    .A2(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6264_ (.A1(_2437_),
    .A2(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6265_ (.A1(_0218_),
    .A2(_3089_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6266_ (.A1(_0211_),
    .A2(\dspArea_regA[21] ),
    .Z(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6267_ (.A1(_0207_),
    .A2(\dspArea_regA[22] ),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6268_ (.A1(_2443_),
    .A2(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6269_ (.A1(_2442_),
    .A2(_2445_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6270_ (.A1(_0213_),
    .A2(_3094_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _6271_ (.A1(_2315_),
    .A2(_2447_),
    .B1(_2382_),
    .B2(_2379_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6272_ (.A1(_2441_),
    .A2(_2446_),
    .A3(_2448_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6273_ (.A1(_2436_),
    .A2(_2449_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6274_ (.A1(_2435_),
    .A2(_2450_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6275_ (.A1(_2432_),
    .A2(_2451_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6276_ (.A1(_2353_),
    .A2(_2362_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6277_ (.A1(_2353_),
    .A2(_2362_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6278_ (.A1(_2453_),
    .A2(_2454_),
    .A3(_2366_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6279_ (.A1(_2367_),
    .A2(_2389_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6280_ (.A1(_2455_),
    .A2(_2456_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6281_ (.A1(_2452_),
    .A2(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6282_ (.A1(_0238_),
    .A2(_3066_),
    .A3(_2401_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6283_ (.A1(_0244_),
    .A2(_3062_),
    .A3(_2403_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6284_ (.A1(_2459_),
    .A2(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6285_ (.I(_2370_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6286_ (.A1(_2373_),
    .A2(_2388_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6287_ (.A1(_2373_),
    .A2(_2388_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6288_ (.A1(_2462_),
    .A2(_2463_),
    .B(_2464_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6289_ (.A1(_0228_),
    .A2(_3081_),
    .A3(_2310_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6290_ (.A1(_0972_),
    .A2(_3070_),
    .A3(_2377_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6291_ (.A1(_2466_),
    .A2(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6292_ (.A1(_0237_),
    .A2(_3070_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6293_ (.A1(_2468_),
    .A2(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6294_ (.A1(_0241_),
    .A2(_3066_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6295_ (.A1(_2470_),
    .A2(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6296_ (.A1(_2465_),
    .A2(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6297_ (.A1(_2461_),
    .A2(_2473_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6298_ (.A1(_2391_),
    .A2(_2394_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6299_ (.A1(_2391_),
    .A2(_2394_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6300_ (.A1(_2475_),
    .A2(_2407_),
    .B(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6301_ (.A1(_2458_),
    .A2(_2474_),
    .A3(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6302_ (.A1(_2399_),
    .A2(_2405_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6303_ (.A1(_2396_),
    .A2(_2406_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6304_ (.A1(_2479_),
    .A2(_2480_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6305_ (.A1(_2478_),
    .A2(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6306_ (.A1(_2408_),
    .A2(_2411_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6307_ (.A1(_2408_),
    .A2(_2411_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6308_ (.A1(_2351_),
    .A2(_2483_),
    .B(_2484_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6309_ (.A1(_2482_),
    .A2(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6310_ (.A1(_2351_),
    .A2(_2483_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6311_ (.A1(_2351_),
    .A2(_2483_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6312_ (.A1(_2348_),
    .A2(_2487_),
    .A3(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6313_ (.A1(_2268_),
    .A2(_2331_),
    .B(_2412_),
    .C(_2347_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6314_ (.A1(_2415_),
    .A2(_2416_),
    .A3(_2333_),
    .A4(_2490_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6315_ (.A1(_2489_),
    .A2(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6316_ (.A1(_2334_),
    .A2(_2413_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6317_ (.I(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6318_ (.A1(_2337_),
    .A2(_2340_),
    .A3(_2343_),
    .B(_2494_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6319_ (.A1(_2492_),
    .A2(_2495_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6320_ (.A1(_2486_),
    .A2(_2496_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6321_ (.I0(\dspArea_regP[30] ),
    .I1(_2497_),
    .S(_0874_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6322_ (.A1(_3111_),
    .A2(_2498_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6323_ (.I(\dspArea_regP[31] ),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6324_ (.I(_2482_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6325_ (.A1(_2500_),
    .A2(_2485_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6326_ (.A1(_2500_),
    .A2(_2485_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6327_ (.A1(_2492_),
    .A2(_2495_),
    .B(_2502_),
    .C(_2501_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6328_ (.A1(_2458_),
    .A2(_2474_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6329_ (.A1(_2458_),
    .A2(_2474_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6330_ (.A1(_2504_),
    .A2(_2505_),
    .A3(_2477_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6331_ (.A1(_2478_),
    .A2(_2481_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6332_ (.A1(\dspArea_regP[30] ),
    .A2(_2428_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6333_ (.I(_0203_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6334_ (.I(_3106_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6335_ (.A1(_2509_),
    .A2(_2510_),
    .A3(_2355_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6336_ (.A1(\dspArea_regP[31] ),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6337_ (.A1(_2508_),
    .A2(_2512_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6338_ (.I(_2441_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6339_ (.A1(_2446_),
    .A2(_2448_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6340_ (.A1(_2446_),
    .A2(_2448_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6341_ (.A1(_2514_),
    .A2(_2515_),
    .B(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6342_ (.A1(_2423_),
    .A2(_2424_),
    .A3(_2427_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6343_ (.A1(_0232_),
    .A2(_3080_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6344_ (.A1(_0227_),
    .A2(_3085_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6345_ (.A1(_0222_),
    .A2(_3089_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6346_ (.A1(_2520_),
    .A2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6347_ (.A1(_2519_),
    .A2(_2522_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6348_ (.A1(_0634_),
    .A2(_3093_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6349_ (.A1(_0211_),
    .A2(_3097_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6350_ (.A1(_0207_),
    .A2(_3101_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6351_ (.A1(_2525_),
    .A2(_2526_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6352_ (.A1(_2524_),
    .A2(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6353_ (.A1(_0207_),
    .A2(_3098_),
    .A3(_2443_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6354_ (.A1(_2442_),
    .A2(_2445_),
    .B(_2529_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6355_ (.A1(_2523_),
    .A2(_2528_),
    .A3(_2530_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6356_ (.A1(_2518_),
    .A2(_2531_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6357_ (.A1(_2517_),
    .A2(_2532_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6358_ (.A1(_2513_),
    .A2(_2533_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6359_ (.A1(_2429_),
    .A2(_2431_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6360_ (.A1(_2432_),
    .A2(_2451_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6361_ (.A1(_2535_),
    .A2(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6362_ (.A1(_2534_),
    .A2(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6363_ (.I(_2468_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6364_ (.A1(_2539_),
    .A2(_2469_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6365_ (.A1(_0243_),
    .A2(_3066_),
    .A3(_2470_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6366_ (.A1(_2540_),
    .A2(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6367_ (.A1(_2436_),
    .A2(_2449_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6368_ (.A1(_2435_),
    .A2(_2450_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6369_ (.A1(_2543_),
    .A2(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6370_ (.A1(_0228_),
    .A2(_3086_),
    .A3(_2376_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6371_ (.A1(_0972_),
    .A2(_3076_),
    .A3(_2440_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6372_ (.A1(_2546_),
    .A2(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6373_ (.A1(_0237_),
    .A2(_3076_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6374_ (.A1(_2548_),
    .A2(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6375_ (.A1(_0241_),
    .A2(_3070_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6376_ (.A1(_2550_),
    .A2(_2551_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6377_ (.A1(_2545_),
    .A2(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6378_ (.A1(_2542_),
    .A2(_2553_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6379_ (.A1(_2538_),
    .A2(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6380_ (.I(_2452_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6381_ (.A1(_2556_),
    .A2(_2457_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6382_ (.A1(_2557_),
    .A2(_2505_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6383_ (.A1(_2465_),
    .A2(_2472_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6384_ (.A1(_2459_),
    .A2(_2460_),
    .B(_2473_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6385_ (.A1(_2559_),
    .A2(_2560_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6386_ (.A1(_2555_),
    .A2(_2558_),
    .A3(_2561_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6387_ (.A1(_2506_),
    .A2(_2507_),
    .A3(_2562_),
    .Z(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6388_ (.A1(_2506_),
    .A2(_2507_),
    .B(_2562_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6389_ (.A1(_2563_),
    .A2(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6390_ (.I(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6391_ (.A1(_2501_),
    .A2(_2503_),
    .A3(_2566_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6392_ (.A1(_2501_),
    .A2(_2503_),
    .B(_2566_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6393_ (.A1(_0792_),
    .A2(_2567_),
    .A3(_2568_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6394_ (.A1(_2499_),
    .A2(_0297_),
    .B(_2569_),
    .C(_1461_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6395_ (.A1(\dspArea_regP[31] ),
    .A2(_2511_),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6396_ (.A1(\dspArea_regP[32] ),
    .A2(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6397_ (.A1(_2421_),
    .A2(_2422_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6398_ (.I(_2523_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6399_ (.A1(_2528_),
    .A2(_2530_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6400_ (.A1(_2528_),
    .A2(_2530_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6401_ (.A1(_2573_),
    .A2(_2574_),
    .B(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6402_ (.A1(_0232_),
    .A2(_3086_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6403_ (.A1(_0227_),
    .A2(_3089_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6404_ (.A1(_0222_),
    .A2(_3093_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6405_ (.A1(_2578_),
    .A2(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6406_ (.A1(_2577_),
    .A2(_2580_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6407_ (.A1(_0211_),
    .A2(_3101_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6408_ (.A1(_0207_),
    .A2(\dspArea_regA[24] ),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6409_ (.A1(_2582_),
    .A2(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6410_ (.A1(_0219_),
    .A2(_3098_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6411_ (.A1(_2584_),
    .A2(_2585_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6412_ (.A1(_0213_),
    .A2(_3102_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6413_ (.A1(_2444_),
    .A2(_2587_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6414_ (.A1(_0219_),
    .A2(_3094_),
    .A3(_2527_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6415_ (.A1(_2588_),
    .A2(_2589_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6416_ (.A1(_2581_),
    .A2(_2586_),
    .A3(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6417_ (.A1(_2572_),
    .A2(_2576_),
    .A3(_2591_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6418_ (.A1(_2571_),
    .A2(_2592_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6419_ (.A1(_2508_),
    .A2(_2512_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6420_ (.A1(_2513_),
    .A2(_2533_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6421_ (.A1(_2594_),
    .A2(_2595_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6422_ (.A1(_2593_),
    .A2(_2596_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6423_ (.I(_2548_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6424_ (.A1(_2598_),
    .A2(_2549_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6425_ (.A1(_2550_),
    .A2(_2551_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6426_ (.A1(_2599_),
    .A2(_2600_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6427_ (.A1(_2518_),
    .A2(_2531_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6428_ (.A1(_2517_),
    .A2(_2532_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6429_ (.A1(_2602_),
    .A2(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6430_ (.A1(_0229_),
    .A2(_3090_),
    .A3(_2439_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6431_ (.A1(_0234_),
    .A2(_3081_),
    .A3(_2522_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6432_ (.A1(_2605_),
    .A2(_2606_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6433_ (.A1(_0238_),
    .A2(_3081_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6434_ (.A1(_2607_),
    .A2(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6435_ (.A1(_0242_),
    .A2(_3076_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6436_ (.A1(_2609_),
    .A2(_2610_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6437_ (.A1(_2604_),
    .A2(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6438_ (.A1(_2601_),
    .A2(_2612_),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6439_ (.A1(_2597_),
    .A2(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6440_ (.I(_2534_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6441_ (.A1(_2615_),
    .A2(_2537_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6442_ (.A1(_2538_),
    .A2(_2554_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6443_ (.A1(_2616_),
    .A2(_2617_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6444_ (.A1(_2614_),
    .A2(_2618_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6445_ (.A1(_2545_),
    .A2(_2552_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6446_ (.A1(_2542_),
    .A2(_2553_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6447_ (.A1(_2620_),
    .A2(_2621_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6448_ (.I(_2622_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6449_ (.A1(_2619_),
    .A2(_2623_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6450_ (.A1(_2555_),
    .A2(_2558_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6451_ (.A1(_2555_),
    .A2(_2558_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6452_ (.A1(_2626_),
    .A2(_2561_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6453_ (.A1(_2625_),
    .A2(_2627_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6454_ (.A1(_2624_),
    .A2(_2628_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _6455_ (.A1(_2624_),
    .A2(_2628_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6456_ (.A1(_2629_),
    .A2(_2630_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6457_ (.A1(_1964_),
    .A2(_2070_),
    .A3(_2161_),
    .A4(_2260_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6458_ (.A1(_2334_),
    .A2(_2413_),
    .A3(_2486_),
    .A4(_2565_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6459_ (.A1(_2632_),
    .A2(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6460_ (.A1(_2489_),
    .A2(_2491_),
    .B(_2565_),
    .C(_2486_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6461_ (.A1(_2501_),
    .A2(_2563_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6462_ (.A1(_2564_),
    .A2(_2635_),
    .A3(_2636_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6463_ (.A1(_2337_),
    .A2(_2340_),
    .B(_2633_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6464_ (.A1(_2634_),
    .A2(_2637_),
    .A3(_2638_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6465_ (.A1(_1967_),
    .A2(_1970_),
    .A3(_2637_),
    .A4(_2638_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6466_ (.A1(_1974_),
    .A2(_2640_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6467_ (.A1(_2639_),
    .A2(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6468_ (.A1(_2631_),
    .A2(_2642_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6469_ (.I0(\dspArea_regP[32] ),
    .I1(_2643_),
    .S(_0874_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6470_ (.A1(_3111_),
    .A2(_2644_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6471_ (.I(\dspArea_regP[33] ),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6472_ (.A1(_2631_),
    .A2(_2642_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6473_ (.A1(_2614_),
    .A2(_2618_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6474_ (.A1(_2619_),
    .A2(_2623_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6475_ (.A1(_2647_),
    .A2(_2648_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6476_ (.A1(_0213_),
    .A2(_3105_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6477_ (.A1(_0634_),
    .A2(_3102_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6478_ (.A1(_2650_),
    .A2(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6479_ (.A1(_2587_),
    .A2(_2583_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6480_ (.A1(_2584_),
    .A2(_2585_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6481_ (.A1(_2653_),
    .A2(_2654_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6482_ (.A1(_2652_),
    .A2(_2655_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6483_ (.A1(_0972_),
    .A2(_3090_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6484_ (.A1(_0227_),
    .A2(_3093_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6485_ (.A1(_0223_),
    .A2(_3097_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6486_ (.A1(_2658_),
    .A2(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6487_ (.A1(_2657_),
    .A2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6488_ (.A1(_2656_),
    .A2(_2661_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6489_ (.A1(_2588_),
    .A2(_2589_),
    .B(_2586_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6490_ (.A1(_2588_),
    .A2(_2589_),
    .A3(_2586_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6491_ (.A1(_2581_),
    .A2(_2664_),
    .A3(_2663_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6492_ (.A1(_2663_),
    .A2(_2665_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6493_ (.A1(_2662_),
    .A2(_2666_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6494_ (.A1(_2645_),
    .A2(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6495_ (.A1(\dspArea_regP[32] ),
    .A2(_2570_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6496_ (.A1(_2571_),
    .A2(_2592_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6497_ (.A1(_2669_),
    .A2(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6498_ (.A1(_2668_),
    .A2(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6499_ (.I(_2607_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6500_ (.A1(_2673_),
    .A2(_2608_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6501_ (.A1(_2609_),
    .A2(_2610_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6502_ (.A1(_2674_),
    .A2(_2675_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6503_ (.A1(_2573_),
    .A2(_2574_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6504_ (.A1(_2575_),
    .A2(_2677_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6505_ (.A1(_2572_),
    .A2(_2591_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6506_ (.A1(_2572_),
    .A2(_2591_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6507_ (.A1(_2678_),
    .A2(_2679_),
    .B(_2680_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6508_ (.A1(_0229_),
    .A2(_3094_),
    .A3(_2521_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6509_ (.A1(_0972_),
    .A2(_3086_),
    .A3(_2580_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6510_ (.A1(_2682_),
    .A2(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6511_ (.A1(_0237_),
    .A2(_3086_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6512_ (.A1(_2684_),
    .A2(_2685_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6513_ (.A1(_0242_),
    .A2(_3081_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6514_ (.A1(_2686_),
    .A2(_2687_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6515_ (.A1(_2681_),
    .A2(_2688_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6516_ (.A1(_2676_),
    .A2(_2689_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6517_ (.A1(_2672_),
    .A2(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6518_ (.I(_2593_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6519_ (.A1(_2692_),
    .A2(_2596_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6520_ (.A1(_2597_),
    .A2(_2613_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6521_ (.A1(_2693_),
    .A2(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6522_ (.A1(_2691_),
    .A2(_2695_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6523_ (.A1(_2604_),
    .A2(_2611_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6524_ (.A1(_2601_),
    .A2(_2612_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6525_ (.A1(_2697_),
    .A2(_2698_),
    .Z(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6526_ (.A1(_2696_),
    .A2(_2699_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6527_ (.A1(_2649_),
    .A2(_2700_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6528_ (.A1(_2630_),
    .A2(_2646_),
    .A3(_2701_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6529_ (.A1(_2630_),
    .A2(_2646_),
    .B(_2701_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6530_ (.A1(_0792_),
    .A2(_2702_),
    .A3(_2703_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6531_ (.A1(_2645_),
    .A2(_0297_),
    .B(_2704_),
    .C(_1461_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6532_ (.A1(\dspArea_regP[33] ),
    .A2(_2667_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6533_ (.A1(_0972_),
    .A2(_3094_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6534_ (.A1(_0227_),
    .A2(_3098_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6535_ (.A1(_0223_),
    .A2(_3102_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6536_ (.A1(_2707_),
    .A2(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6537_ (.A1(_2706_),
    .A2(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6538_ (.A1(_0219_),
    .A2(_3106_),
    .A3(_2582_),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6539_ (.A1(_2710_),
    .A2(_2711_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6540_ (.I(_2655_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6541_ (.A1(_2652_),
    .A2(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6542_ (.A1(_2656_),
    .A2(_2661_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6543_ (.A1(_2714_),
    .A2(_2715_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6544_ (.A1(_2712_),
    .A2(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6545_ (.A1(\dspArea_regP[34] ),
    .A2(_2717_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6546_ (.A1(_2705_),
    .A2(_2718_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6547_ (.I(_2684_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6548_ (.A1(_2720_),
    .A2(_2685_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6549_ (.A1(_2686_),
    .A2(_2687_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6550_ (.A1(_2721_),
    .A2(_2722_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6551_ (.I(_2662_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6552_ (.A1(_2724_),
    .A2(_2666_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6553_ (.A1(_0229_),
    .A2(_3098_),
    .A3(_2579_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6554_ (.A1(_0234_),
    .A2(_3090_),
    .A3(_2660_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6555_ (.A1(_2726_),
    .A2(_2727_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6556_ (.A1(_0237_),
    .A2(_3090_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6557_ (.A1(_2728_),
    .A2(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6558_ (.A1(_0242_),
    .A2(_3086_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6559_ (.A1(_2730_),
    .A2(_2731_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6560_ (.A1(_2725_),
    .A2(_2732_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6561_ (.A1(_2723_),
    .A2(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6562_ (.A1(_2719_),
    .A2(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6563_ (.I(_2671_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6564_ (.A1(_2668_),
    .A2(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6565_ (.A1(_2672_),
    .A2(_2690_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6566_ (.A1(_2737_),
    .A2(_2738_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6567_ (.A1(_2735_),
    .A2(_2739_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6568_ (.A1(_2681_),
    .A2(_2688_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6569_ (.A1(_2676_),
    .A2(_2689_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6570_ (.A1(_2741_),
    .A2(_2742_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6571_ (.A1(_2740_),
    .A2(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6572_ (.A1(_2691_),
    .A2(_2695_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6573_ (.A1(_2696_),
    .A2(_2699_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6574_ (.A1(_2745_),
    .A2(_2746_),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6575_ (.A1(_2744_),
    .A2(_2747_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6576_ (.A1(_2649_),
    .A2(_2700_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6577_ (.A1(_2649_),
    .A2(_2700_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6578_ (.A1(_2630_),
    .A2(_2750_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6579_ (.A1(_2629_),
    .A2(_2630_),
    .A3(_2701_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6580_ (.I(_2752_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6581_ (.A1(_1974_),
    .A2(_2640_),
    .B(_2753_),
    .C(_2639_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6582_ (.A1(_2749_),
    .A2(_2751_),
    .A3(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6583_ (.A1(_2748_),
    .A2(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6584_ (.I0(\dspArea_regP[34] ),
    .I1(_2756_),
    .S(_0874_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6585_ (.A1(_3111_),
    .A2(_2757_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6586_ (.I(\dspArea_regP[35] ),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6587_ (.A1(_2735_),
    .A2(_2739_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6588_ (.A1(_2740_),
    .A2(_2743_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6589_ (.A1(\dspArea_regP[34] ),
    .A2(_2717_),
    .Z(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6590_ (.A1(_0234_),
    .A2(_3098_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6591_ (.A1(_0228_),
    .A2(_3102_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6592_ (.A1(_0223_),
    .A2(_3105_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6593_ (.A1(_2763_),
    .A2(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6594_ (.A1(_2762_),
    .A2(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6595_ (.A1(_2587_),
    .A2(_2710_),
    .B(_0219_),
    .C(_3106_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6596_ (.A1(_2766_),
    .A2(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6597_ (.A1(_2758_),
    .A2(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6598_ (.A1(_2761_),
    .A2(_2769_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6599_ (.I(_2728_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6600_ (.A1(_2771_),
    .A2(_2729_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6601_ (.A1(_2730_),
    .A2(_2731_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6602_ (.A1(_2772_),
    .A2(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6603_ (.I(_2712_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6604_ (.A1(_2775_),
    .A2(_2716_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6605_ (.A1(_2659_),
    .A2(_2763_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6606_ (.A1(_0234_),
    .A2(_3094_),
    .A3(_2709_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6607_ (.A1(_0238_),
    .A2(_3094_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6608_ (.A1(_2777_),
    .A2(_2778_),
    .A3(_2779_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6609_ (.A1(_2777_),
    .A2(_2778_),
    .B(_2779_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6610_ (.A1(_2780_),
    .A2(_2781_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6611_ (.A1(_0243_),
    .A2(_3090_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6612_ (.A1(_2782_),
    .A2(_2783_),
    .Z(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6613_ (.A1(_2776_),
    .A2(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6614_ (.A1(_2774_),
    .A2(_2785_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6615_ (.A1(_2770_),
    .A2(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6616_ (.A1(_2705_),
    .A2(_2718_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6617_ (.A1(_2719_),
    .A2(_2734_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6618_ (.A1(_2788_),
    .A2(_2789_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6619_ (.A1(_2725_),
    .A2(_2732_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6620_ (.A1(_2723_),
    .A2(_2733_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6621_ (.A1(_2791_),
    .A2(_2792_),
    .Z(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _6622_ (.A1(_2787_),
    .A2(_2790_),
    .A3(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6623_ (.A1(_2759_),
    .A2(_2760_),
    .A3(_2794_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6624_ (.A1(_2759_),
    .A2(_2760_),
    .B(_2794_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6625_ (.A1(_2795_),
    .A2(_2796_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6626_ (.I(_2748_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6627_ (.A1(_2744_),
    .A2(_2747_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6628_ (.A1(_2798_),
    .A2(_2755_),
    .B(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6629_ (.A1(_2797_),
    .A2(_2800_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6630_ (.A1(_0792_),
    .A2(_2801_),
    .Z(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6631_ (.A1(_2758_),
    .A2(_0297_),
    .B(_2802_),
    .C(_1461_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6632_ (.A1(_2748_),
    .A2(_2752_),
    .A3(_2797_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6633_ (.A1(_1974_),
    .A2(_2640_),
    .B(_2803_),
    .C(_2639_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6634_ (.A1(_2630_),
    .A2(_2749_),
    .B(_2750_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6635_ (.A1(_2748_),
    .A2(_2797_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6636_ (.I(_2795_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6637_ (.A1(_2799_),
    .A2(_2807_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6638_ (.A1(_2805_),
    .A2(_2806_),
    .B(_2808_),
    .C(_2796_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6639_ (.A1(\dspArea_regP[35] ),
    .A2(_2768_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6640_ (.A1(_0229_),
    .A2(_3106_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6641_ (.A1(_0234_),
    .A2(_3102_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6642_ (.A1(_2811_),
    .A2(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6643_ (.A1(\dspArea_regP[36] ),
    .A2(_2813_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6644_ (.A1(_2810_),
    .A2(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6645_ (.A1(_2782_),
    .A2(_2783_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6646_ (.A1(_2781_),
    .A2(_2816_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6647_ (.I(_2767_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6648_ (.A1(_2766_),
    .A2(_2818_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6649_ (.A1(_0223_),
    .A2(_3106_),
    .A3(_2763_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6650_ (.A1(_0234_),
    .A2(_3098_),
    .A3(_2765_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6651_ (.A1(_0238_),
    .A2(_3098_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6652_ (.A1(_2820_),
    .A2(_2821_),
    .A3(_2822_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6653_ (.A1(_2820_),
    .A2(_2821_),
    .B(_2822_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6654_ (.A1(_2823_),
    .A2(_2824_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6655_ (.A1(_0243_),
    .A2(_3094_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6656_ (.A1(_2825_),
    .A2(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6657_ (.A1(_2819_),
    .A2(_2827_),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6658_ (.A1(_2817_),
    .A2(_2828_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6659_ (.A1(_2815_),
    .A2(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6660_ (.A1(_2761_),
    .A2(_2769_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6661_ (.A1(_2770_),
    .A2(_2786_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6662_ (.A1(_2831_),
    .A2(_2832_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6663_ (.A1(_2830_),
    .A2(_2833_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6664_ (.A1(_2776_),
    .A2(_2784_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6665_ (.A1(_2774_),
    .A2(_2785_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6666_ (.A1(_2835_),
    .A2(_2836_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6667_ (.A1(_2834_),
    .A2(_2837_),
    .Z(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6668_ (.A1(_2787_),
    .A2(_2790_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6669_ (.A1(_2787_),
    .A2(_2790_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6670_ (.A1(_2840_),
    .A2(_2793_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6671_ (.A1(_2839_),
    .A2(_2841_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6672_ (.A1(_2838_),
    .A2(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6673_ (.A1(_2804_),
    .A2(_2809_),
    .B(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6674_ (.A1(_2843_),
    .A2(_2804_),
    .A3(_2809_),
    .Z(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6675_ (.A1(_2844_),
    .A2(_2845_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6676_ (.A1(\dspArea_regP[36] ),
    .A2(_0874_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6677_ (.A1(_0299_),
    .A2(_2846_),
    .B(_2847_),
    .C(_1461_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6678_ (.A1(\dspArea_regP[37] ),
    .A2(_0259_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6679_ (.I(_2838_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6680_ (.A1(_2849_),
    .A2(_2842_),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6681_ (.A1(_2850_),
    .A2(_2844_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6682_ (.I(_2833_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6683_ (.A1(_2830_),
    .A2(_2852_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6684_ (.A1(_2834_),
    .A2(_2837_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6685_ (.A1(\dspArea_regP[36] ),
    .A2(_2813_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6686_ (.A1(_0234_),
    .A2(_3106_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6687_ (.A1(\dspArea_regP[37] ),
    .A2(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6688_ (.A1(_2855_),
    .A2(_2857_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6689_ (.A1(_0238_),
    .A2(_3102_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6690_ (.A1(_2763_),
    .A2(_2856_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6691_ (.I0(_2859_),
    .I1(_0238_),
    .S(_2860_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6692_ (.A1(_0243_),
    .A2(_3098_),
    .Z(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6693_ (.A1(_2861_),
    .A2(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6694_ (.A1(_0244_),
    .A2(_3094_),
    .A3(_2825_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6695_ (.A1(_2824_),
    .A2(_2864_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6696_ (.A1(_2863_),
    .A2(_2865_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6697_ (.A1(_2858_),
    .A2(_2866_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6698_ (.A1(_2810_),
    .A2(_2814_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6699_ (.I(_2815_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6700_ (.A1(_2869_),
    .A2(_2829_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6701_ (.A1(_2868_),
    .A2(_2870_),
    .Z(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6702_ (.A1(_2867_),
    .A2(_2871_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6703_ (.A1(_2819_),
    .A2(_2827_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6704_ (.I(_2817_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6705_ (.A1(_2874_),
    .A2(_2828_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6706_ (.A1(_2873_),
    .A2(_2875_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6707_ (.A1(_2872_),
    .A2(_2876_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6708_ (.A1(_2853_),
    .A2(_2854_),
    .A3(_2877_),
    .Z(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6709_ (.A1(_2853_),
    .A2(_2854_),
    .B(_2877_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6710_ (.A1(_2878_),
    .A2(_2879_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6711_ (.A1(_2851_),
    .A2(_2880_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6712_ (.A1(_0259_),
    .A2(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6713_ (.A1(_3110_),
    .A2(_2848_),
    .A3(_2882_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6714_ (.I(_2865_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6715_ (.A1(_2863_),
    .A2(_2883_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6716_ (.A1(\dspArea_regP[37] ),
    .A2(_2856_),
    .Z(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6717_ (.A1(\dspArea_regP[38] ),
    .A2(_2885_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6718_ (.A1(_0238_),
    .A2(_3106_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6719_ (.A1(_0243_),
    .A2(_3102_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6720_ (.A1(_2887_),
    .A2(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6721_ (.A1(_0238_),
    .A2(_2860_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6722_ (.I(_2861_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6723_ (.A1(_2891_),
    .A2(_2862_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6724_ (.A1(_2890_),
    .A2(_2892_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6725_ (.A1(_2889_),
    .A2(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6726_ (.A1(_2886_),
    .A2(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6727_ (.A1(_2855_),
    .A2(_2857_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6728_ (.A1(_2858_),
    .A2(_2866_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6729_ (.A1(_2896_),
    .A2(_2897_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6730_ (.A1(_2895_),
    .A2(_2898_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6731_ (.A1(_2884_),
    .A2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6732_ (.A1(_2867_),
    .A2(_2871_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6733_ (.A1(_2872_),
    .A2(_2876_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6734_ (.A1(_2901_),
    .A2(_2902_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6735_ (.A1(_2900_),
    .A2(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6736_ (.A1(_2850_),
    .A2(_2879_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6737_ (.A1(_2844_),
    .A2(_2905_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6738_ (.A1(_2878_),
    .A2(_2906_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6739_ (.A1(_2904_),
    .A2(_2907_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6740_ (.A1(\dspArea_regP[38] ),
    .A2(_0299_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6741_ (.A1(_0299_),
    .A2(_2908_),
    .B(_2909_),
    .C(_3109_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6742_ (.I(\dspArea_regP[39] ),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6743_ (.A1(_2900_),
    .A2(_2903_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6744_ (.I(_2878_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6745_ (.A1(_2844_),
    .A2(_2905_),
    .B(_2904_),
    .C(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6746_ (.A1(_2889_),
    .A2(_2893_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6747_ (.A1(_0244_),
    .A2(_3106_),
    .A3(_2859_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6748_ (.A1(\dspArea_regP[39] ),
    .A2(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6749_ (.A1(\dspArea_regP[38] ),
    .A2(_2885_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6750_ (.A1(_2886_),
    .A2(_2894_),
    .Z(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6751_ (.A1(_2917_),
    .A2(_2918_),
    .Z(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6752_ (.A1(_2916_),
    .A2(_2919_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6753_ (.A1(_2914_),
    .A2(_2920_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6754_ (.A1(_2884_),
    .A2(_2899_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6755_ (.A1(_2895_),
    .A2(_2898_),
    .B(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6756_ (.A1(_2921_),
    .A2(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6757_ (.A1(_2921_),
    .A2(_2923_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6758_ (.A1(_2924_),
    .A2(_2925_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6759_ (.A1(_2911_),
    .A2(_2913_),
    .B(_2926_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6760_ (.A1(_2911_),
    .A2(_2913_),
    .A3(_2926_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6761_ (.A1(_0874_),
    .A2(_2927_),
    .A3(_2928_),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6762_ (.A1(_2910_),
    .A2(_0297_),
    .B(_2929_),
    .C(_3109_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6763_ (.A1(_2904_),
    .A2(_2926_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6764_ (.A1(_2843_),
    .A2(_2880_),
    .A3(_2930_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6765_ (.A1(_2809_),
    .A2(_2931_),
    .Z(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6766_ (.A1(_2878_),
    .A2(_2930_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6767_ (.A1(_2911_),
    .A2(_2925_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6768_ (.A1(_2905_),
    .A2(_2933_),
    .B1(_2934_),
    .B2(_2924_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6769_ (.A1(_2804_),
    .A2(_2931_),
    .B(_2932_),
    .C(_2935_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6770_ (.A1(_2916_),
    .A2(_2919_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6771_ (.A1(_2914_),
    .A2(_2920_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6772_ (.A1(_2937_),
    .A2(_2938_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6773_ (.I(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6774_ (.I(_0244_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6775_ (.A1(_2910_),
    .A2(_2859_),
    .B(_2510_),
    .C(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6776_ (.A1(\dspArea_regP[40] ),
    .A2(_2942_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6777_ (.A1(_2940_),
    .A2(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6778_ (.A1(_2936_),
    .A2(_2944_),
    .Z(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6779_ (.I0(\dspArea_regP[40] ),
    .I1(_2945_),
    .S(_0874_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6780_ (.A1(_3111_),
    .A2(_2946_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6781_ (.A1(\dspArea_regP[40] ),
    .A2(_2942_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6782_ (.A1(\dspArea_regP[41] ),
    .A2(_2947_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6783_ (.A1(\dspArea_regP[41] ),
    .A2(_2947_),
    .Z(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6784_ (.A1(_2948_),
    .A2(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6785_ (.A1(_2940_),
    .A2(_2943_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6786_ (.A1(_2936_),
    .A2(_2944_),
    .B(_2951_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6787_ (.A1(_2950_),
    .A2(_2952_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6788_ (.A1(\dspArea_regP[41] ),
    .A2(_0874_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6789_ (.A1(_0792_),
    .A2(_2953_),
    .B(_2954_),
    .C(_3109_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _6790_ (.A1(_2944_),
    .A2(_2950_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6791_ (.A1(_2951_),
    .A2(_2948_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6792_ (.A1(_2949_),
    .A2(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6793_ (.A1(_2936_),
    .A2(_2955_),
    .B(_2957_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6794_ (.A1(_0298_),
    .A2(_2958_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6795_ (.A1(\dspArea_regP[42] ),
    .A2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _6796_ (.A1(\dspArea_regP[42] ),
    .A2(_0250_),
    .A3(_2958_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6797_ (.A1(_3142_),
    .A2(_2960_),
    .A3(_2961_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6798_ (.A1(\dspArea_regP[43] ),
    .A2(_2961_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6799_ (.A1(_3111_),
    .A2(_2962_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6800_ (.A1(\dspArea_regP[43] ),
    .A2(\dspArea_regP[42] ),
    .Z(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6801_ (.I(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6802_ (.A1(\dspArea_regP[43] ),
    .A2(\dspArea_regP[42] ),
    .A3(_2949_),
    .A4(_2956_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6803_ (.A1(_2936_),
    .A2(_2955_),
    .A3(_2964_),
    .B(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6804_ (.A1(_0250_),
    .A2(_2966_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _6805_ (.A1(\dspArea_regP[44] ),
    .A2(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6806_ (.A1(_3112_),
    .A2(_2968_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6807_ (.A1(\dspArea_regP[44] ),
    .A2(_0298_),
    .A3(_2958_),
    .A4(_2963_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6808_ (.A1(\dspArea_regP[45] ),
    .A2(_2969_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6809_ (.A1(\dspArea_regP[45] ),
    .A2(\dspArea_regP[44] ),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6810_ (.A1(_0298_),
    .A2(_2958_),
    .A3(_2963_),
    .A4(_2971_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6811_ (.A1(_3142_),
    .A2(_2970_),
    .A3(_2972_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6812_ (.A1(\dspArea_regP[46] ),
    .A2(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6813_ (.A1(\dspArea_regP[46] ),
    .A2(_0250_),
    .A3(_2966_),
    .A4(_2971_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6814_ (.A1(_3142_),
    .A2(_2973_),
    .A3(_2974_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6815_ (.A1(\dspArea_regP[47] ),
    .A2(_2974_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6816_ (.A1(_3111_),
    .A2(_2975_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6817_ (.D(_0125_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(_zz_1_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6818_ (.D(_0126_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6819_ (.D(_0127_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6820_ (.D(_0128_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6821_ (.D(_0129_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6822_ (.D(_0130_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6823_ (.D(_0131_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6824_ (.D(_0132_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6825_ (.D(_0133_),
    .CLK(net65),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6826_ (.D(_0134_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6827_ (.D(_0135_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6828_ (.D(_0136_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6829_ (.D(_0137_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6830_ (.D(_0138_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6831_ (.D(_0139_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6832_ (.D(_0140_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6833_ (.D(_0141_),
    .CLK(net65),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6834_ (.D(_0142_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6835_ (.D(_0143_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6836_ (.D(_0144_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6837_ (.D(_0145_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6838_ (.D(_0146_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6839_ (.D(_0147_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6840_ (.D(_0148_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6841_ (.D(_0149_),
    .CLK(net65),
    .Q(net145));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6842_ (.D(_0150_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6843_ (.D(_0151_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6844_ (.D(_0152_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6845_ (.D(_0153_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6846_ (.D(_0000_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6847_ (.D(_0001_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6848_ (.D(_0002_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6849_ (.D(_0003_),
    .CLK(net65),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6850_ (.D(_0004_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6851_ (.D(_0005_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6852_ (.D(_0006_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6853_ (.D(_0007_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6854_ (.D(_0008_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6855_ (.D(_0009_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6856_ (.D(_0010_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6857_ (.D(_0011_),
    .CLK(net65),
    .Q(net147));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6858_ (.D(_0012_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6859_ (.D(_0013_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6860_ (.D(_0014_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6861_ (.D(_0015_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6862_ (.D(_0016_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6863_ (.D(_0017_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6864_ (.D(_0018_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6865_ (.D(_0019_),
    .CLK(net65),
    .Q(net148));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6866_ (.D(_0020_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6867_ (.D(_0021_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6868_ (.D(_0022_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6869_ (.D(_0023_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6870_ (.D(_0024_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6871_ (.D(_0025_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6872_ (.D(_0026_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6873_ (.D(_0027_),
    .CLK(net65),
    .Q(net150));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6874_ (.D(_0028_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6875_ (.D(_0029_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6876_ (.D(_0030_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6877_ (.D(_0031_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6878_ (.D(_0032_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6879_ (.D(_0033_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6880_ (.D(_0034_),
    .CLK(net65),
    .Q(\dacArea_dac_cnt_7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6881_ (.D(_0035_),
    .CLK(net65),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6882_ (.D(_0036_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6883_ (.D(_0037_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6884_ (.D(_0038_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6885_ (.D(_0039_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6886_ (.D(_0040_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6887_ (.D(_0041_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6888_ (.D(_0042_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6889_ (.D(_0043_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6890_ (.D(_0044_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6891_ (.D(_0045_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6892_ (.D(_0046_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6893_ (.D(_0047_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6894_ (.D(_0048_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regA[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6895_ (.D(_0049_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6896_ (.D(_0050_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6897_ (.D(_0051_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6898_ (.D(_0052_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regA[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6899_ (.D(_0053_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regA[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6900_ (.D(_0054_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regA[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6901_ (.D(_0055_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regA[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6902_ (.D(_0056_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6903_ (.D(_0057_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6904_ (.D(_0058_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6905_ (.D(_0059_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6906_ (.D(_0060_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6907_ (.D(_0061_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6908_ (.D(_0062_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6909_ (.D(_0063_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6910_ (.D(_0064_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6911_ (.D(_0065_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6912_ (.D(_0066_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6913_ (.D(_0067_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6914_ (.D(_0068_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6915_ (.D(_0069_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6916_ (.D(_0070_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6917_ (.D(_0071_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6918_ (.D(_0072_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regB[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6919_ (.D(_0073_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\dspArea_regB[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6920_ (.D(_0074_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6921_ (.D(_0075_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regB[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6922_ (.D(_0076_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regB[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6923_ (.D(_0077_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6924_ (.D(_0078_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6925_ (.D(_0079_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6926_ (.D(_0080_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6927_ (.D(_0081_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6928_ (.D(_0082_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6929_ (.D(_0083_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6930_ (.D(_0084_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6931_ (.D(_0085_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6932_ (.D(_0086_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6933_ (.D(_0087_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6934_ (.D(_0088_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6935_ (.D(_0089_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6936_ (.D(_0090_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6937_ (.D(_0091_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6938_ (.D(_0092_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6939_ (.D(_0093_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6940_ (.D(_0094_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6941_ (.D(_0095_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6942_ (.D(_0096_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6943_ (.D(_0097_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6944_ (.D(_0098_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6945_ (.D(_0099_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6946_ (.D(_0100_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6947_ (.D(_0101_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6948_ (.D(_0102_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6949_ (.D(_0103_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6950_ (.D(_0104_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6951_ (.D(_0105_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6952_ (.D(_0106_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6953_ (.D(_0107_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6954_ (.D(_0108_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6955_ (.D(_0109_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6956_ (.D(_0110_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6957_ (.D(_0111_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6958_ (.D(_0112_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6959_ (.D(_0113_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6960_ (.D(_0114_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6961_ (.D(_0115_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6962_ (.D(_0116_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6963_ (.D(_0117_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6964_ (.D(_0118_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6965_ (.D(_0119_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6966_ (.D(_0120_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6967_ (.D(_0121_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6968_ (.D(_0122_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6969_ (.D(_0123_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6970_ (.D(_0124_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\dspArea_regP[47] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_199 (.Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_200 (.Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_201 (.Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_202 (.Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_203 (.Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_204 (.Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_205 (.Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_206 (.Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_207 (.Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_208 (.Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_209 (.Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_210 (.Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_211 (.Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_212 (.Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_213 (.Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_214 (.Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_215 (.Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_216 (.Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_217 (.Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_218 (.Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_219 (.Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_220 (.Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_221 (.Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_222 (.Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_223 (.Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_224 (.Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_225 (.Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_226 (.Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_227 (.Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_228 (.Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_229 (.Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_230 (.Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_231 (.Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_232 (.Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_233 (.Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_234 (.Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_235 (.Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tieh DSP48_198 (.Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7015_ (.I(net143),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7016_ (.I(net144),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7017_ (.I(net145),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7018_ (.I(net146),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(net147),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7020_ (.I(net148),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7021_ (.I(net150),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7022_ (.I(net151),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7023_ (.I(net143),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7024_ (.I(net144),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7025_ (.I(net145),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7026_ (.I(net146),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7027_ (.I(net147),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7028_ (.I(net148),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7029_ (.I(net150),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7030_ (.I(net151),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7031_ (.I(net143),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7032_ (.I(net144),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7033_ (.I(net145),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7034_ (.I(net146),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7035_ (.I(net147),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7036_ (.I(net148),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7037_ (.I(net150),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7038_ (.I(net151),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(la_data_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(la_data_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(la_data_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(la_data_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(la_data_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(la_data_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(la_data_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(la_data_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(la_data_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(la_data_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(la_data_in[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(la_data_in[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(la_data_in[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(la_data_in[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(la_data_in[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(la_data_in[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(la_data_in[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(la_data_in[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(la_data_in[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(la_data_in[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(la_data_in[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(la_data_in[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(la_data_in[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(la_data_in[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(la_data_in[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(la_data_in[32]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(la_data_in[33]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(la_data_in[34]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(la_data_in[35]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input30 (.I(la_data_in[36]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input31 (.I(la_data_in[37]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input32 (.I(la_data_in[38]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(la_data_in[39]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(la_data_in[3]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(la_data_in[40]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(la_data_in[41]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input37 (.I(la_data_in[42]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input38 (.I(la_data_in[43]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(la_data_in[44]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(la_data_in[45]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(la_data_in[46]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(la_data_in[47]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(la_data_in[48]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(la_data_in[49]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input45 (.I(la_data_in[4]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(la_data_in[50]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(la_data_in[51]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(la_data_in[52]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(la_data_in[53]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input50 (.I(la_data_in[54]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(la_data_in[55]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(la_data_in[56]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(la_data_in[57]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input54 (.I(la_data_in[58]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input55 (.I(la_data_in[59]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input56 (.I(la_data_in[5]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input57 (.I(la_data_in[60]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input58 (.I(la_data_in[61]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input59 (.I(la_data_in[62]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(la_data_in[63]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input61 (.I(la_data_in[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(la_data_in[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(la_data_in[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(la_data_in[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 input65 (.I(user_clock2),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(wb_ADR[0]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(wb_ADR[10]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(wb_ADR[11]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(wb_ADR[12]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(wb_ADR[13]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(wb_ADR[14]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(wb_ADR[15]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(wb_ADR[16]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(wb_ADR[17]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(wb_ADR[18]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(wb_ADR[19]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(wb_ADR[1]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(wb_ADR[20]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(wb_ADR[21]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(wb_ADR[22]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(wb_ADR[23]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input82 (.I(wb_ADR[24]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input83 (.I(wb_ADR[25]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input84 (.I(wb_ADR[26]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(wb_ADR[27]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(wb_ADR[28]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(wb_ADR[29]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(wb_ADR[2]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(wb_ADR[30]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input90 (.I(wb_ADR[31]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input91 (.I(wb_ADR[3]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input92 (.I(wb_ADR[4]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input93 (.I(wb_ADR[5]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input94 (.I(wb_ADR[6]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input95 (.I(wb_ADR[7]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input96 (.I(wb_ADR[8]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input97 (.I(wb_ADR[9]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input98 (.I(wb_CYC),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input99 (.I(wb_DAT_MOSI[0]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input100 (.I(wb_DAT_MOSI[10]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input101 (.I(wb_DAT_MOSI[11]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input102 (.I(wb_DAT_MOSI[12]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input103 (.I(wb_DAT_MOSI[13]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input104 (.I(wb_DAT_MOSI[14]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input105 (.I(wb_DAT_MOSI[15]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input106 (.I(wb_DAT_MOSI[16]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input107 (.I(wb_DAT_MOSI[17]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input108 (.I(wb_DAT_MOSI[18]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input109 (.I(wb_DAT_MOSI[19]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input110 (.I(wb_DAT_MOSI[1]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input111 (.I(wb_DAT_MOSI[20]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input112 (.I(wb_DAT_MOSI[21]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input113 (.I(wb_DAT_MOSI[22]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input114 (.I(wb_DAT_MOSI[23]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input115 (.I(wb_DAT_MOSI[24]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input116 (.I(wb_DAT_MOSI[2]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input117 (.I(wb_DAT_MOSI[3]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input118 (.I(wb_DAT_MOSI[4]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input119 (.I(wb_DAT_MOSI[5]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input120 (.I(wb_DAT_MOSI[6]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input121 (.I(wb_DAT_MOSI[7]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input122 (.I(wb_DAT_MOSI[8]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input123 (.I(wb_DAT_MOSI[9]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input124 (.I(wb_STB),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input125 (.I(wb_WE),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input126 (.I(wb_rst_i),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output127 (.I(net127),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output128 (.I(net128),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output129 (.I(net129),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output130 (.I(net130),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output131 (.I(net131),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output132 (.I(net132),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output133 (.I(net133),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output134 (.I(net134),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output135 (.I(net135),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output136 (.I(net136),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output137 (.I(net137),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output138 (.I(net138),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output139 (.I(net139),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output140 (.I(net140),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output141 (.I(net141),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output142 (.I(net142),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output143 (.I(net143),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output144 (.I(net144),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output145 (.I(net145),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output146 (.I(net146),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output147 (.I(net147),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output148 (.I(net148),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output149 (.I(net149),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output150 (.I(net150),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output151 (.I(net151),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output152 (.I(net152),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output153 (.I(net153),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output154 (.I(net154),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output155 (.I(net155),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output156 (.I(net156),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output157 (.I(net157),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output158 (.I(net158),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output159 (.I(net159),
    .Z(wb_ACK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output160 (.I(net160),
    .Z(wb_DAT_MISO[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output161 (.I(net161),
    .Z(wb_DAT_MISO[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output162 (.I(net162),
    .Z(wb_DAT_MISO[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output163 (.I(net163),
    .Z(wb_DAT_MISO[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output164 (.I(net164),
    .Z(wb_DAT_MISO[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output165 (.I(net165),
    .Z(wb_DAT_MISO[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output166 (.I(net166),
    .Z(wb_DAT_MISO[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output167 (.I(net167),
    .Z(wb_DAT_MISO[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output168 (.I(net168),
    .Z(wb_DAT_MISO[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output169 (.I(net169),
    .Z(wb_DAT_MISO[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output170 (.I(net170),
    .Z(wb_DAT_MISO[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output171 (.I(net171),
    .Z(wb_DAT_MISO[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output172 (.I(net172),
    .Z(wb_DAT_MISO[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output173 (.I(net173),
    .Z(wb_DAT_MISO[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output174 (.I(net174),
    .Z(wb_DAT_MISO[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output175 (.I(net175),
    .Z(wb_DAT_MISO[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output176 (.I(net176),
    .Z(wb_DAT_MISO[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output177 (.I(net177),
    .Z(wb_DAT_MISO[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output178 (.I(net178),
    .Z(wb_DAT_MISO[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output179 (.I(net179),
    .Z(wb_DAT_MISO[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output180 (.I(net180),
    .Z(wb_DAT_MISO[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output181 (.I(net181),
    .Z(wb_DAT_MISO[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output182 (.I(net182),
    .Z(wb_DAT_MISO[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output183 (.I(net183),
    .Z(wb_DAT_MISO[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output184 (.I(net184),
    .Z(wb_DAT_MISO[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output185 (.I(net185),
    .Z(wb_DAT_MISO[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output186 (.I(net186),
    .Z(wb_DAT_MISO[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output187 (.I(net187),
    .Z(wb_DAT_MISO[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output188 (.I(net188),
    .Z(wb_DAT_MISO[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output189 (.I(net189),
    .Z(wb_DAT_MISO[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output190 (.I(net190),
    .Z(wb_DAT_MISO[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output191 (.I(net191),
    .Z(wb_DAT_MISO[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSP48_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__D (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__D (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__D (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A1 (.I(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__C (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A1 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I0 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__S (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__S (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__I (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__I (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I0 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__I0 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__I (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__I (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__I (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I0 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__I (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__I (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__I0 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__I0 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__I (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__I (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__I0 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__I (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__I (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__I (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__I0 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__I (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__I (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__I0 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__I (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__I (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__I0 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__I (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__I (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__I (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__B (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I0 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__I (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__I (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I0 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__I (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__I (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__I (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__I (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__I0 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__I (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__I (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__I (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__I0 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__I (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__I1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__I0 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__I (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__I (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__I (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__I (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I0 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A3 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__I (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__B (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A3 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__S (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__S (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__S (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__S (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__I (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__I (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__B (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A3 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A3 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A3 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__I1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__S (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__I (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A3 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A3 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__I (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__I1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A3 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A3 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A3 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A3 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A3 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A3 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A3 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__I (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A3 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__C (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A3 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__S (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__S (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__S (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__S (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A3 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A3 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A3 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A3 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A3 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A3 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__I (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A3 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A3 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A3 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__B (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A3 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__B (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A3 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A3 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__B (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A3 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__I (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A3 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A1 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A3 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__B (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A3 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__B (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__C (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__C (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A3 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A3 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A3 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A2 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A3 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__B (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A3 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__C (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__I (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A3 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A3 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A3 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__B (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__B (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A2 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A3 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A3 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__B (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A3 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A3 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__I (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A3 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__B (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A3 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A3 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A3 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A3 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__B (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A3 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A3 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__B (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A3 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A3 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__B (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__B (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__I1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__I (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A3 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A3 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__I (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A3 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A3 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__B (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A3 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A3 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__I (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A3 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__B (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A3 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A3 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__I (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__I (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A3 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A3 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__B (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__I (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A3 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A4 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__B1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__C (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__I (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A3 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A3 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A3 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A3 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A3 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A3 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A3 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A3 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A3 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__B (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A3 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__C (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__I (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A3 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A3 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A3 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__B (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__I (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A3 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__B (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A3 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__B (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A3 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A3 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__I1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A2 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A3 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A3 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A3 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A3 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__I1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__B (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__I (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A3 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__B (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A3 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A4 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__I (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__B (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A2 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A2 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A2 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A3 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A4 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A3 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__C (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__C (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__I (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__I1 (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A3 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A3 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A1 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__B (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A2 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A3 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__I (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A3 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A3 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A1 (.I(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A3 (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__I (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__B1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__B1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__B1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__B1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__B1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__I (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__I (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__B1 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__I (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__I (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A3 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__B2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__I (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__C1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__C1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__I (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__C1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__C1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__C1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__C1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__I (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__B2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__I (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__I (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__I (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__B2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__I (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__I (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__B2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__I (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__I (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__C1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__I (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__I (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A3 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__I (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__B2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__I (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__I (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__I (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__B2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__I (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__I (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A4 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__B2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__I (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__I (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A4 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A3 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__B2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__I (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A4 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A3 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__I (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__B2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__I (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A3 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__I (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__B2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__I (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__I (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__I (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__B2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__I (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__I (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__B2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__I (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__I (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__B2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__I (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__I (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__I (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__B2 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__I (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__I (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__I (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__B2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__I (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__I (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__I (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__I (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__I (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__I (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__I (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__I (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__I (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A1 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__I (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__I (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A1 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__I (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A3 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__I (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__C (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__I (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__C (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__C (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__C (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A3 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A1 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A4 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A3 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A1 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A2 (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A2 (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__I (.I(\dspArea_regA[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__I (.I(\dspArea_regA[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A2 (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I (.I(\dspArea_regA[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A2 (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A3 (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__I (.I(\dspArea_regA[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(\dspArea_regB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(\dspArea_regB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__I (.I(\dspArea_regB[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__I (.I(\dspArea_regB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__C2 (.I(\dspArea_regP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I0 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__C2 (.I(\dspArea_regP[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__C2 (.I(\dspArea_regP[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I0 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__C2 (.I(\dspArea_regP[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__C2 (.I(\dspArea_regP[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__C2 (.I(\dspArea_regP[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__C2 (.I(\dspArea_regP[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I0 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(\dspArea_regP[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A1 (.I(\dspArea_regP[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I0 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A1 (.I(\dspArea_regP[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(\dspArea_regP[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(\dspArea_regP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__I0 (.I(\dspArea_regP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(\dspArea_regP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__C2 (.I(\dspArea_regP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I0 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A1 (.I(\dspArea_regP[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__I (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(\dspArea_regP[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__I0 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(\dspArea_regP[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A1 (.I(\dspArea_regP[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I0 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A1 (.I(\dspArea_regP[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__I (.I(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(\dspArea_regP[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A1 (.I(\dspArea_regP[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__I0 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(\dspArea_regP[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A1 (.I(\dspArea_regP[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__I0 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__C2 (.I(\dspArea_regP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__I0 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(\dspArea_regP[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__I (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A1 (.I(\dspArea_regP[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__I0 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A1 (.I(\dspArea_regP[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__I (.I(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(\dspArea_regP[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__I0 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A1 (.I(\dspArea_regP[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A1 (.I(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__I (.I(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A1 (.I(\dspArea_regP[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(\dspArea_regP[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(\dspArea_regP[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A1 (.I(\dspArea_regP[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__I (.I(\dspArea_regP[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(\dspArea_regP[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__I0 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__C2 (.I(\dspArea_regP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A1 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__I0 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A1 (.I(\dspArea_regP[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A1 (.I(\dspArea_regP[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A2 (.I(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A2 (.I(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A1 (.I(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A1 (.I(\dspArea_regP[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(\dspArea_regP[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A2 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__A1 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A1 (.I(\dspArea_regP[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A1 (.I(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A1 (.I(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(\dspArea_regP[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A1 (.I(\dspArea_regP[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A1 (.I(\dspArea_regP[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(\dspArea_regP[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__I (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__C2 (.I(\dspArea_regP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__C2 (.I(\dspArea_regP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__I0 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__C2 (.I(\dspArea_regP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__I0 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__C2 (.I(\dspArea_regP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A1 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__C2 (.I(\dspArea_regP[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__I0 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__C2 (.I(\dspArea_regP[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(la_data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(la_data_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(la_data_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(la_data_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(la_data_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(la_data_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(la_data_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(la_data_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(la_data_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(la_data_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(la_data_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(la_data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(la_data_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(la_data_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(la_data_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(la_data_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(la_data_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(la_data_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(la_data_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(la_data_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(la_data_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(la_data_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(la_data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(la_data_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(la_data_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(la_data_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(la_data_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(la_data_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(la_data_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(la_data_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(la_data_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(la_data_in[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(la_data_in[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(la_data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(la_data_in[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(la_data_in[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(la_data_in[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(la_data_in[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(la_data_in[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(la_data_in[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(la_data_in[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(la_data_in[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(la_data_in[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(la_data_in[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(la_data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(la_data_in[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(la_data_in[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(la_data_in[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(la_data_in[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(la_data_in[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(la_data_in[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(la_data_in[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(la_data_in[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(la_data_in[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(la_data_in[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(la_data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(la_data_in[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(la_data_in[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(la_data_in[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(la_data_in[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(la_data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(la_data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(la_data_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(la_data_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(user_clock2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(wb_ADR[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(wb_ADR[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(wb_ADR[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(wb_ADR[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(wb_ADR[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(wb_ADR[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(wb_ADR[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(wb_ADR[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(wb_ADR[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(wb_ADR[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(wb_ADR[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(wb_ADR[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(wb_ADR[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(wb_ADR[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(wb_ADR[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(wb_ADR[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(wb_ADR[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(wb_ADR[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(wb_ADR[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(wb_ADR[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(wb_ADR[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(wb_ADR[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(wb_ADR[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(wb_ADR[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(wb_ADR[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(wb_ADR[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(wb_ADR[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(wb_ADR[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(wb_ADR[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(wb_ADR[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(wb_ADR[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(wb_ADR[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(wb_CYC));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(wb_DAT_MOSI[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(wb_DAT_MOSI[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(wb_DAT_MOSI[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(wb_DAT_MOSI[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(wb_DAT_MOSI[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(wb_DAT_MOSI[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(wb_DAT_MOSI[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(wb_DAT_MOSI[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(wb_DAT_MOSI[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(wb_DAT_MOSI[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(wb_DAT_MOSI[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(wb_DAT_MOSI[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(wb_DAT_MOSI[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(wb_DAT_MOSI[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(wb_DAT_MOSI[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(wb_DAT_MOSI[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(wb_DAT_MOSI[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(wb_DAT_MOSI[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(wb_DAT_MOSI[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(wb_DAT_MOSI[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(wb_DAT_MOSI[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(wb_DAT_MOSI[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(wb_DAT_MOSI[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(wb_DAT_MOSI[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(wb_DAT_MOSI[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(wb_STB));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(wb_WE));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A2 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A3 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__I1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__I1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__I1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__I1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__I1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__I1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__I1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__I1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__I1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__I1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A2 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A1 (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output144_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output146_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output167_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net198;
 assign io_oeb[10] = net208;
 assign io_oeb[11] = net209;
 assign io_oeb[12] = net210;
 assign io_oeb[13] = net211;
 assign io_oeb[14] = net212;
 assign io_oeb[15] = net213;
 assign io_oeb[16] = net214;
 assign io_oeb[17] = net215;
 assign io_oeb[18] = net216;
 assign io_oeb[19] = net217;
 assign io_oeb[1] = net199;
 assign io_oeb[20] = net218;
 assign io_oeb[21] = net219;
 assign io_oeb[22] = net220;
 assign io_oeb[23] = net221;
 assign io_oeb[24] = net222;
 assign io_oeb[25] = net223;
 assign io_oeb[26] = net224;
 assign io_oeb[27] = net225;
 assign io_oeb[28] = net226;
 assign io_oeb[29] = net227;
 assign io_oeb[2] = net200;
 assign io_oeb[30] = net228;
 assign io_oeb[31] = net229;
 assign io_oeb[32] = net230;
 assign io_oeb[33] = net231;
 assign io_oeb[34] = net232;
 assign io_oeb[35] = net233;
 assign io_oeb[36] = net234;
 assign io_oeb[37] = net235;
 assign io_oeb[3] = net201;
 assign io_oeb[4] = net202;
 assign io_oeb[5] = net203;
 assign io_oeb[6] = net204;
 assign io_oeb[7] = net205;
 assign io_oeb[8] = net206;
 assign io_oeb[9] = net207;
 assign io_out[32] = net192;
 assign io_out[33] = net193;
 assign io_out[34] = net194;
 assign io_out[35] = net195;
 assign io_out[36] = net196;
 assign io_out[37] = net197;
endmodule

