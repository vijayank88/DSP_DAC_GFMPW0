VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSP48
  CLASS BLOCK ;
  FOREIGN DSP48 ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 596.000 7.280 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 596.000 242.480 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 596.000 266.000 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 596.000 289.520 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 596.000 313.040 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 596.000 336.560 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 596.000 360.080 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 596.000 383.600 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 596.000 407.120 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 596.000 430.640 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 596.000 454.160 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 596.000 30.800 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 596.000 477.680 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 596.000 501.200 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 596.000 524.720 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 596.000 548.240 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 596.000 571.760 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 596.000 595.280 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 596.000 618.800 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 596.000 642.320 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 596.000 665.840 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 596.000 689.360 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 596.000 54.320 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 596.000 712.880 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 596.000 736.400 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 596.000 759.920 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 596.000 783.440 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 596.000 806.960 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 596.000 830.480 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 596.000 854.000 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 596.000 877.520 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 596.000 77.840 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 596.000 101.360 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 596.000 124.880 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 596.000 148.400 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 596.000 171.920 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 596.000 195.440 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 596.000 218.960 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 596.000 15.120 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 596.000 250.320 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 596.000 273.840 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 596.000 297.360 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 596.000 320.880 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 596.000 344.400 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 596.000 367.920 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 596.000 391.440 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 596.000 414.960 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 596.000 438.480 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 596.000 462.000 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 596.000 38.640 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 596.000 485.520 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 596.000 509.040 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 596.000 532.560 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 596.000 556.080 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 596.000 579.600 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 596.000 603.120 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 626.080 596.000 626.640 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 596.000 650.160 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.120 596.000 673.680 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 596.000 697.200 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 596.000 62.160 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 596.000 720.720 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 596.000 744.240 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 596.000 767.760 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 596.000 791.280 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.240 596.000 814.800 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 596.000 838.320 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 596.000 861.840 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 596.000 885.360 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 596.000 85.680 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 596.000 109.200 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 596.000 132.720 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 596.000 156.240 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 596.000 179.760 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 596.000 203.280 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 596.000 226.800 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 596.000 22.960 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 596.000 258.160 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 596.000 281.680 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 596.000 305.200 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 596.000 328.720 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 596.000 352.240 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 596.000 375.760 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 596.000 399.280 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 596.000 422.800 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 596.000 446.320 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 596.000 469.840 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 596.000 46.480 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.800 596.000 493.360 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 596.000 516.880 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 596.000 540.400 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.360 596.000 563.920 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.880 596.000 587.440 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 596.000 610.960 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 596.000 634.480 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 657.440 596.000 658.000 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 596.000 681.520 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 596.000 705.040 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 596.000 70.000 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 596.000 728.560 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 596.000 752.080 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 775.040 596.000 775.600 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 798.560 596.000 799.120 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 596.000 822.640 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 845.600 596.000 846.160 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 869.120 596.000 869.680 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 596.000 893.200 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 596.000 93.520 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 596.000 117.040 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 596.000 140.560 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 596.000 164.080 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 596.000 187.600 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 596.000 211.120 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 596.000 234.640 600.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 0.000 598.640 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 603.120 0.000 603.680 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 0.000 608.720 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 613.200 0.000 613.760 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 0.000 618.800 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 623.280 0.000 623.840 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 0.000 628.880 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.360 0.000 633.920 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 0.000 638.960 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 643.440 0.000 644.000 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.720 0.000 553.280 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 0.000 649.040 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 653.520 0.000 654.080 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 0.000 659.120 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 663.600 0.000 664.160 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 0.000 669.200 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 673.680 0.000 674.240 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 683.760 0.000 684.320 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 0.000 689.360 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.840 0.000 694.400 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 0.000 558.320 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 0.000 699.440 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 703.920 0.000 704.480 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 0.000 709.520 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.000 0.000 714.560 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 0.000 719.600 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 724.080 0.000 724.640 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 0.000 729.680 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 734.160 0.000 734.720 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 0.000 739.760 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 744.240 0.000 744.800 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 562.800 0.000 563.360 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 754.320 0.000 754.880 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 0.000 759.920 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 764.400 0.000 764.960 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 0.000 770.000 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 774.480 0.000 775.040 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 0.000 780.080 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 784.560 0.000 785.120 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 0.000 790.160 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.640 0.000 795.200 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 0.000 568.400 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 0.000 800.240 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 804.720 0.000 805.280 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 0.000 810.320 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 814.800 0.000 815.360 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 0.000 820.400 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 824.880 0.000 825.440 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 0.000 830.480 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 834.960 0.000 835.520 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 0.000 840.560 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 845.040 0.000 845.600 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 572.880 0.000 573.440 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 0.000 850.640 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 855.120 0.000 855.680 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 0.000 860.720 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 865.200 0.000 865.760 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 0.000 578.480 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 582.960 0.000 583.520 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 593.040 0.000 593.600 4.000 ;
    END
  END la_data_in[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 0.000 870.800 4.000 ;
    END
  END user_clock2
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 584.380 ;
    END
  END vss
  PIN wb_ACK
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.560 0.000 29.120 4.000 ;
    END
  END wb_ACK
  PIN wb_ADR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END wb_ADR[0]
  PIN wb_ADR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END wb_ADR[10]
  PIN wb_ADR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.160 0.000 230.720 4.000 ;
    END
  END wb_ADR[11]
  PIN wb_ADR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 0.000 245.840 4.000 ;
    END
  END wb_ADR[12]
  PIN wb_ADR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.400 0.000 260.960 4.000 ;
    END
  END wb_ADR[13]
  PIN wb_ADR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END wb_ADR[14]
  PIN wb_ADR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.640 0.000 291.200 4.000 ;
    END
  END wb_ADR[15]
  PIN wb_ADR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END wb_ADR[16]
  PIN wb_ADR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.880 0.000 321.440 4.000 ;
    END
  END wb_ADR[17]
  PIN wb_ADR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 0.000 336.560 4.000 ;
    END
  END wb_ADR[18]
  PIN wb_ADR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.120 0.000 351.680 4.000 ;
    END
  END wb_ADR[19]
  PIN wb_ADR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.960 0.000 79.520 4.000 ;
    END
  END wb_ADR[1]
  PIN wb_ADR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 0.000 366.800 4.000 ;
    END
  END wb_ADR[20]
  PIN wb_ADR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.360 0.000 381.920 4.000 ;
    END
  END wb_ADR[21]
  PIN wb_ADR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END wb_ADR[22]
  PIN wb_ADR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.600 0.000 412.160 4.000 ;
    END
  END wb_ADR[23]
  PIN wb_ADR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END wb_ADR[24]
  PIN wb_ADR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.840 0.000 442.400 4.000 ;
    END
  END wb_ADR[25]
  PIN wb_ADR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 0.000 457.520 4.000 ;
    END
  END wb_ADR[26]
  PIN wb_ADR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.080 0.000 472.640 4.000 ;
    END
  END wb_ADR[27]
  PIN wb_ADR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 0.000 487.760 4.000 ;
    END
  END wb_ADR[28]
  PIN wb_ADR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 502.320 0.000 502.880 4.000 ;
    END
  END wb_ADR[29]
  PIN wb_ADR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END wb_ADR[2]
  PIN wb_ADR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END wb_ADR[30]
  PIN wb_ADR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.560 0.000 533.120 4.000 ;
    END
  END wb_ADR[31]
  PIN wb_ADR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.200 0.000 109.760 4.000 ;
    END
  END wb_ADR[3]
  PIN wb_ADR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END wb_ADR[4]
  PIN wb_ADR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 139.440 0.000 140.000 4.000 ;
    END
  END wb_ADR[5]
  PIN wb_ADR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END wb_ADR[6]
  PIN wb_ADR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.680 0.000 170.240 4.000 ;
    END
  END wb_ADR[7]
  PIN wb_ADR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END wb_ADR[8]
  PIN wb_ADR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.920 0.000 200.480 4.000 ;
    END
  END wb_ADR[9]
  PIN wb_CYC
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END wb_CYC
  PIN wb_DAT_MISO[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.880 0.000 69.440 4.000 ;
    END
  END wb_DAT_MISO[0]
  PIN wb_DAT_MISO[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.080 0.000 220.640 4.000 ;
    END
  END wb_DAT_MISO[10]
  PIN wb_DAT_MISO[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END wb_DAT_MISO[11]
  PIN wb_DAT_MISO[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 250.320 0.000 250.880 4.000 ;
    END
  END wb_DAT_MISO[12]
  PIN wb_DAT_MISO[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END wb_DAT_MISO[13]
  PIN wb_DAT_MISO[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.560 0.000 281.120 4.000 ;
    END
  END wb_DAT_MISO[14]
  PIN wb_DAT_MISO[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 0.000 296.240 4.000 ;
    END
  END wb_DAT_MISO[15]
  PIN wb_DAT_MISO[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.800 0.000 311.360 4.000 ;
    END
  END wb_DAT_MISO[16]
  PIN wb_DAT_MISO[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 0.000 326.480 4.000 ;
    END
  END wb_DAT_MISO[17]
  PIN wb_DAT_MISO[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.040 0.000 341.600 4.000 ;
    END
  END wb_DAT_MISO[18]
  PIN wb_DAT_MISO[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END wb_DAT_MISO[19]
  PIN wb_DAT_MISO[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END wb_DAT_MISO[1]
  PIN wb_DAT_MISO[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.280 0.000 371.840 4.000 ;
    END
  END wb_DAT_MISO[20]
  PIN wb_DAT_MISO[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END wb_DAT_MISO[21]
  PIN wb_DAT_MISO[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 401.520 0.000 402.080 4.000 ;
    END
  END wb_DAT_MISO[22]
  PIN wb_DAT_MISO[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 0.000 417.200 4.000 ;
    END
  END wb_DAT_MISO[23]
  PIN wb_DAT_MISO[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.760 0.000 432.320 4.000 ;
    END
  END wb_DAT_MISO[24]
  PIN wb_DAT_MISO[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 0.000 447.440 4.000 ;
    END
  END wb_DAT_MISO[25]
  PIN wb_DAT_MISO[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.000 0.000 462.560 4.000 ;
    END
  END wb_DAT_MISO[26]
  PIN wb_DAT_MISO[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 0.000 477.680 4.000 ;
    END
  END wb_DAT_MISO[27]
  PIN wb_DAT_MISO[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.240 0.000 492.800 4.000 ;
    END
  END wb_DAT_MISO[28]
  PIN wb_DAT_MISO[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END wb_DAT_MISO[29]
  PIN wb_DAT_MISO[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.120 0.000 99.680 4.000 ;
    END
  END wb_DAT_MISO[2]
  PIN wb_DAT_MISO[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 522.480 0.000 523.040 4.000 ;
    END
  END wb_DAT_MISO[30]
  PIN wb_DAT_MISO[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 0.000 538.160 4.000 ;
    END
  END wb_DAT_MISO[31]
  PIN wb_DAT_MISO[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END wb_DAT_MISO[3]
  PIN wb_DAT_MISO[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.360 0.000 129.920 4.000 ;
    END
  END wb_DAT_MISO[4]
  PIN wb_DAT_MISO[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END wb_DAT_MISO[5]
  PIN wb_DAT_MISO[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.600 0.000 160.160 4.000 ;
    END
  END wb_DAT_MISO[6]
  PIN wb_DAT_MISO[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END wb_DAT_MISO[7]
  PIN wb_DAT_MISO[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.840 0.000 190.400 4.000 ;
    END
  END wb_DAT_MISO[8]
  PIN wb_DAT_MISO[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END wb_DAT_MISO[9]
  PIN wb_DAT_MOSI[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END wb_DAT_MOSI[0]
  PIN wb_DAT_MOSI[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END wb_DAT_MOSI[10]
  PIN wb_DAT_MOSI[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 240.240 0.000 240.800 4.000 ;
    END
  END wb_DAT_MOSI[11]
  PIN wb_DAT_MOSI[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END wb_DAT_MOSI[12]
  PIN wb_DAT_MOSI[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.480 0.000 271.040 4.000 ;
    END
  END wb_DAT_MOSI[13]
  PIN wb_DAT_MOSI[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 0.000 286.160 4.000 ;
    END
  END wb_DAT_MOSI[14]
  PIN wb_DAT_MOSI[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.720 0.000 301.280 4.000 ;
    END
  END wb_DAT_MOSI[15]
  PIN wb_DAT_MOSI[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END wb_DAT_MOSI[16]
  PIN wb_DAT_MOSI[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.960 0.000 331.520 4.000 ;
    END
  END wb_DAT_MOSI[17]
  PIN wb_DAT_MOSI[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END wb_DAT_MOSI[18]
  PIN wb_DAT_MOSI[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 361.200 0.000 361.760 4.000 ;
    END
  END wb_DAT_MOSI[19]
  PIN wb_DAT_MOSI[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.040 0.000 89.600 4.000 ;
    END
  END wb_DAT_MOSI[1]
  PIN wb_DAT_MOSI[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 0.000 376.880 4.000 ;
    END
  END wb_DAT_MOSI[20]
  PIN wb_DAT_MOSI[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 391.440 0.000 392.000 4.000 ;
    END
  END wb_DAT_MOSI[21]
  PIN wb_DAT_MOSI[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 0.000 407.120 4.000 ;
    END
  END wb_DAT_MOSI[22]
  PIN wb_DAT_MOSI[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.680 0.000 422.240 4.000 ;
    END
  END wb_DAT_MOSI[23]
  PIN wb_DAT_MOSI[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 0.000 437.360 4.000 ;
    END
  END wb_DAT_MOSI[24]
  PIN wb_DAT_MOSI[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.920 0.000 452.480 4.000 ;
    END
  END wb_DAT_MOSI[25]
  PIN wb_DAT_MOSI[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 0.000 467.600 4.000 ;
    END
  END wb_DAT_MOSI[26]
  PIN wb_DAT_MOSI[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 482.160 0.000 482.720 4.000 ;
    END
  END wb_DAT_MOSI[27]
  PIN wb_DAT_MOSI[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 0.000 497.840 4.000 ;
    END
  END wb_DAT_MOSI[28]
  PIN wb_DAT_MOSI[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.400 0.000 512.960 4.000 ;
    END
  END wb_DAT_MOSI[29]
  PIN wb_DAT_MOSI[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END wb_DAT_MOSI[2]
  PIN wb_DAT_MOSI[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 0.000 528.080 4.000 ;
    END
  END wb_DAT_MOSI[30]
  PIN wb_DAT_MOSI[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.640 0.000 543.200 4.000 ;
    END
  END wb_DAT_MOSI[31]
  PIN wb_DAT_MOSI[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.280 0.000 119.840 4.000 ;
    END
  END wb_DAT_MOSI[3]
  PIN wb_DAT_MOSI[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END wb_DAT_MOSI[4]
  PIN wb_DAT_MOSI[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.520 0.000 150.080 4.000 ;
    END
  END wb_DAT_MOSI[5]
  PIN wb_DAT_MOSI[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END wb_DAT_MOSI[6]
  PIN wb_DAT_MOSI[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.760 0.000 180.320 4.000 ;
    END
  END wb_DAT_MOSI[7]
  PIN wb_DAT_MOSI[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END wb_DAT_MOSI[8]
  PIN wb_DAT_MOSI[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.000 0.000 210.560 4.000 ;
    END
  END wb_DAT_MOSI[9]
  PIN wb_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.640 0.000 39.200 4.000 ;
    END
  END wb_SEL
  PIN wb_STB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END wb_STB
  PIN wb_WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 48.720 0.000 49.280 4.000 ;
    END
  END wb_WE
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 0.000 59.360 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 893.200 585.050 ;
      LAYER Metal2 ;
        RECT 7.980 595.700 14.260 596.000 ;
        RECT 15.420 595.700 22.100 596.000 ;
        RECT 23.260 595.700 29.940 596.000 ;
        RECT 31.100 595.700 37.780 596.000 ;
        RECT 38.940 595.700 45.620 596.000 ;
        RECT 46.780 595.700 53.460 596.000 ;
        RECT 54.620 595.700 61.300 596.000 ;
        RECT 62.460 595.700 69.140 596.000 ;
        RECT 70.300 595.700 76.980 596.000 ;
        RECT 78.140 595.700 84.820 596.000 ;
        RECT 85.980 595.700 92.660 596.000 ;
        RECT 93.820 595.700 100.500 596.000 ;
        RECT 101.660 595.700 108.340 596.000 ;
        RECT 109.500 595.700 116.180 596.000 ;
        RECT 117.340 595.700 124.020 596.000 ;
        RECT 125.180 595.700 131.860 596.000 ;
        RECT 133.020 595.700 139.700 596.000 ;
        RECT 140.860 595.700 147.540 596.000 ;
        RECT 148.700 595.700 155.380 596.000 ;
        RECT 156.540 595.700 163.220 596.000 ;
        RECT 164.380 595.700 171.060 596.000 ;
        RECT 172.220 595.700 178.900 596.000 ;
        RECT 180.060 595.700 186.740 596.000 ;
        RECT 187.900 595.700 194.580 596.000 ;
        RECT 195.740 595.700 202.420 596.000 ;
        RECT 203.580 595.700 210.260 596.000 ;
        RECT 211.420 595.700 218.100 596.000 ;
        RECT 219.260 595.700 225.940 596.000 ;
        RECT 227.100 595.700 233.780 596.000 ;
        RECT 234.940 595.700 241.620 596.000 ;
        RECT 242.780 595.700 249.460 596.000 ;
        RECT 250.620 595.700 257.300 596.000 ;
        RECT 258.460 595.700 265.140 596.000 ;
        RECT 266.300 595.700 272.980 596.000 ;
        RECT 274.140 595.700 280.820 596.000 ;
        RECT 281.980 595.700 288.660 596.000 ;
        RECT 289.820 595.700 296.500 596.000 ;
        RECT 297.660 595.700 304.340 596.000 ;
        RECT 305.500 595.700 312.180 596.000 ;
        RECT 313.340 595.700 320.020 596.000 ;
        RECT 321.180 595.700 327.860 596.000 ;
        RECT 329.020 595.700 335.700 596.000 ;
        RECT 336.860 595.700 343.540 596.000 ;
        RECT 344.700 595.700 351.380 596.000 ;
        RECT 352.540 595.700 359.220 596.000 ;
        RECT 360.380 595.700 367.060 596.000 ;
        RECT 368.220 595.700 374.900 596.000 ;
        RECT 376.060 595.700 382.740 596.000 ;
        RECT 383.900 595.700 390.580 596.000 ;
        RECT 391.740 595.700 398.420 596.000 ;
        RECT 399.580 595.700 406.260 596.000 ;
        RECT 407.420 595.700 414.100 596.000 ;
        RECT 415.260 595.700 421.940 596.000 ;
        RECT 423.100 595.700 429.780 596.000 ;
        RECT 430.940 595.700 437.620 596.000 ;
        RECT 438.780 595.700 445.460 596.000 ;
        RECT 446.620 595.700 453.300 596.000 ;
        RECT 454.460 595.700 461.140 596.000 ;
        RECT 462.300 595.700 468.980 596.000 ;
        RECT 470.140 595.700 476.820 596.000 ;
        RECT 477.980 595.700 484.660 596.000 ;
        RECT 485.820 595.700 492.500 596.000 ;
        RECT 493.660 595.700 500.340 596.000 ;
        RECT 501.500 595.700 508.180 596.000 ;
        RECT 509.340 595.700 516.020 596.000 ;
        RECT 517.180 595.700 523.860 596.000 ;
        RECT 525.020 595.700 531.700 596.000 ;
        RECT 532.860 595.700 539.540 596.000 ;
        RECT 540.700 595.700 547.380 596.000 ;
        RECT 548.540 595.700 555.220 596.000 ;
        RECT 556.380 595.700 563.060 596.000 ;
        RECT 564.220 595.700 570.900 596.000 ;
        RECT 572.060 595.700 578.740 596.000 ;
        RECT 579.900 595.700 586.580 596.000 ;
        RECT 587.740 595.700 594.420 596.000 ;
        RECT 595.580 595.700 602.260 596.000 ;
        RECT 603.420 595.700 610.100 596.000 ;
        RECT 611.260 595.700 617.940 596.000 ;
        RECT 619.100 595.700 625.780 596.000 ;
        RECT 626.940 595.700 633.620 596.000 ;
        RECT 634.780 595.700 641.460 596.000 ;
        RECT 642.620 595.700 649.300 596.000 ;
        RECT 650.460 595.700 657.140 596.000 ;
        RECT 658.300 595.700 664.980 596.000 ;
        RECT 666.140 595.700 672.820 596.000 ;
        RECT 673.980 595.700 680.660 596.000 ;
        RECT 681.820 595.700 688.500 596.000 ;
        RECT 689.660 595.700 696.340 596.000 ;
        RECT 697.500 595.700 704.180 596.000 ;
        RECT 705.340 595.700 712.020 596.000 ;
        RECT 713.180 595.700 719.860 596.000 ;
        RECT 721.020 595.700 727.700 596.000 ;
        RECT 728.860 595.700 735.540 596.000 ;
        RECT 736.700 595.700 743.380 596.000 ;
        RECT 744.540 595.700 751.220 596.000 ;
        RECT 752.380 595.700 759.060 596.000 ;
        RECT 760.220 595.700 766.900 596.000 ;
        RECT 768.060 595.700 774.740 596.000 ;
        RECT 775.900 595.700 782.580 596.000 ;
        RECT 783.740 595.700 790.420 596.000 ;
        RECT 791.580 595.700 798.260 596.000 ;
        RECT 799.420 595.700 806.100 596.000 ;
        RECT 807.260 595.700 813.940 596.000 ;
        RECT 815.100 595.700 821.780 596.000 ;
        RECT 822.940 595.700 829.620 596.000 ;
        RECT 830.780 595.700 837.460 596.000 ;
        RECT 838.620 595.700 845.300 596.000 ;
        RECT 846.460 595.700 853.140 596.000 ;
        RECT 854.300 595.700 860.980 596.000 ;
        RECT 862.140 595.700 868.820 596.000 ;
        RECT 869.980 595.700 876.660 596.000 ;
        RECT 877.820 595.700 884.500 596.000 ;
        RECT 885.660 595.700 892.340 596.000 ;
        RECT 7.980 4.300 893.060 595.700 ;
        RECT 7.980 3.500 28.260 4.300 ;
        RECT 29.420 3.500 33.300 4.300 ;
        RECT 34.460 3.500 38.340 4.300 ;
        RECT 39.500 3.500 43.380 4.300 ;
        RECT 44.540 3.500 48.420 4.300 ;
        RECT 49.580 3.500 53.460 4.300 ;
        RECT 54.620 3.500 58.500 4.300 ;
        RECT 59.660 3.500 63.540 4.300 ;
        RECT 64.700 3.500 68.580 4.300 ;
        RECT 69.740 3.500 73.620 4.300 ;
        RECT 74.780 3.500 78.660 4.300 ;
        RECT 79.820 3.500 83.700 4.300 ;
        RECT 84.860 3.500 88.740 4.300 ;
        RECT 89.900 3.500 93.780 4.300 ;
        RECT 94.940 3.500 98.820 4.300 ;
        RECT 99.980 3.500 103.860 4.300 ;
        RECT 105.020 3.500 108.900 4.300 ;
        RECT 110.060 3.500 113.940 4.300 ;
        RECT 115.100 3.500 118.980 4.300 ;
        RECT 120.140 3.500 124.020 4.300 ;
        RECT 125.180 3.500 129.060 4.300 ;
        RECT 130.220 3.500 134.100 4.300 ;
        RECT 135.260 3.500 139.140 4.300 ;
        RECT 140.300 3.500 144.180 4.300 ;
        RECT 145.340 3.500 149.220 4.300 ;
        RECT 150.380 3.500 154.260 4.300 ;
        RECT 155.420 3.500 159.300 4.300 ;
        RECT 160.460 3.500 164.340 4.300 ;
        RECT 165.500 3.500 169.380 4.300 ;
        RECT 170.540 3.500 174.420 4.300 ;
        RECT 175.580 3.500 179.460 4.300 ;
        RECT 180.620 3.500 184.500 4.300 ;
        RECT 185.660 3.500 189.540 4.300 ;
        RECT 190.700 3.500 194.580 4.300 ;
        RECT 195.740 3.500 199.620 4.300 ;
        RECT 200.780 3.500 204.660 4.300 ;
        RECT 205.820 3.500 209.700 4.300 ;
        RECT 210.860 3.500 214.740 4.300 ;
        RECT 215.900 3.500 219.780 4.300 ;
        RECT 220.940 3.500 224.820 4.300 ;
        RECT 225.980 3.500 229.860 4.300 ;
        RECT 231.020 3.500 234.900 4.300 ;
        RECT 236.060 3.500 239.940 4.300 ;
        RECT 241.100 3.500 244.980 4.300 ;
        RECT 246.140 3.500 250.020 4.300 ;
        RECT 251.180 3.500 255.060 4.300 ;
        RECT 256.220 3.500 260.100 4.300 ;
        RECT 261.260 3.500 265.140 4.300 ;
        RECT 266.300 3.500 270.180 4.300 ;
        RECT 271.340 3.500 275.220 4.300 ;
        RECT 276.380 3.500 280.260 4.300 ;
        RECT 281.420 3.500 285.300 4.300 ;
        RECT 286.460 3.500 290.340 4.300 ;
        RECT 291.500 3.500 295.380 4.300 ;
        RECT 296.540 3.500 300.420 4.300 ;
        RECT 301.580 3.500 305.460 4.300 ;
        RECT 306.620 3.500 310.500 4.300 ;
        RECT 311.660 3.500 315.540 4.300 ;
        RECT 316.700 3.500 320.580 4.300 ;
        RECT 321.740 3.500 325.620 4.300 ;
        RECT 326.780 3.500 330.660 4.300 ;
        RECT 331.820 3.500 335.700 4.300 ;
        RECT 336.860 3.500 340.740 4.300 ;
        RECT 341.900 3.500 345.780 4.300 ;
        RECT 346.940 3.500 350.820 4.300 ;
        RECT 351.980 3.500 355.860 4.300 ;
        RECT 357.020 3.500 360.900 4.300 ;
        RECT 362.060 3.500 365.940 4.300 ;
        RECT 367.100 3.500 370.980 4.300 ;
        RECT 372.140 3.500 376.020 4.300 ;
        RECT 377.180 3.500 381.060 4.300 ;
        RECT 382.220 3.500 386.100 4.300 ;
        RECT 387.260 3.500 391.140 4.300 ;
        RECT 392.300 3.500 396.180 4.300 ;
        RECT 397.340 3.500 401.220 4.300 ;
        RECT 402.380 3.500 406.260 4.300 ;
        RECT 407.420 3.500 411.300 4.300 ;
        RECT 412.460 3.500 416.340 4.300 ;
        RECT 417.500 3.500 421.380 4.300 ;
        RECT 422.540 3.500 426.420 4.300 ;
        RECT 427.580 3.500 431.460 4.300 ;
        RECT 432.620 3.500 436.500 4.300 ;
        RECT 437.660 3.500 441.540 4.300 ;
        RECT 442.700 3.500 446.580 4.300 ;
        RECT 447.740 3.500 451.620 4.300 ;
        RECT 452.780 3.500 456.660 4.300 ;
        RECT 457.820 3.500 461.700 4.300 ;
        RECT 462.860 3.500 466.740 4.300 ;
        RECT 467.900 3.500 471.780 4.300 ;
        RECT 472.940 3.500 476.820 4.300 ;
        RECT 477.980 3.500 481.860 4.300 ;
        RECT 483.020 3.500 486.900 4.300 ;
        RECT 488.060 3.500 491.940 4.300 ;
        RECT 493.100 3.500 496.980 4.300 ;
        RECT 498.140 3.500 502.020 4.300 ;
        RECT 503.180 3.500 507.060 4.300 ;
        RECT 508.220 3.500 512.100 4.300 ;
        RECT 513.260 3.500 517.140 4.300 ;
        RECT 518.300 3.500 522.180 4.300 ;
        RECT 523.340 3.500 527.220 4.300 ;
        RECT 528.380 3.500 532.260 4.300 ;
        RECT 533.420 3.500 537.300 4.300 ;
        RECT 538.460 3.500 542.340 4.300 ;
        RECT 543.500 3.500 547.380 4.300 ;
        RECT 548.540 3.500 552.420 4.300 ;
        RECT 553.580 3.500 557.460 4.300 ;
        RECT 558.620 3.500 562.500 4.300 ;
        RECT 563.660 3.500 567.540 4.300 ;
        RECT 568.700 3.500 572.580 4.300 ;
        RECT 573.740 3.500 577.620 4.300 ;
        RECT 578.780 3.500 582.660 4.300 ;
        RECT 583.820 3.500 587.700 4.300 ;
        RECT 588.860 3.500 592.740 4.300 ;
        RECT 593.900 3.500 597.780 4.300 ;
        RECT 598.940 3.500 602.820 4.300 ;
        RECT 603.980 3.500 607.860 4.300 ;
        RECT 609.020 3.500 612.900 4.300 ;
        RECT 614.060 3.500 617.940 4.300 ;
        RECT 619.100 3.500 622.980 4.300 ;
        RECT 624.140 3.500 628.020 4.300 ;
        RECT 629.180 3.500 633.060 4.300 ;
        RECT 634.220 3.500 638.100 4.300 ;
        RECT 639.260 3.500 643.140 4.300 ;
        RECT 644.300 3.500 648.180 4.300 ;
        RECT 649.340 3.500 653.220 4.300 ;
        RECT 654.380 3.500 658.260 4.300 ;
        RECT 659.420 3.500 663.300 4.300 ;
        RECT 664.460 3.500 668.340 4.300 ;
        RECT 669.500 3.500 673.380 4.300 ;
        RECT 674.540 3.500 678.420 4.300 ;
        RECT 679.580 3.500 683.460 4.300 ;
        RECT 684.620 3.500 688.500 4.300 ;
        RECT 689.660 3.500 693.540 4.300 ;
        RECT 694.700 3.500 698.580 4.300 ;
        RECT 699.740 3.500 703.620 4.300 ;
        RECT 704.780 3.500 708.660 4.300 ;
        RECT 709.820 3.500 713.700 4.300 ;
        RECT 714.860 3.500 718.740 4.300 ;
        RECT 719.900 3.500 723.780 4.300 ;
        RECT 724.940 3.500 728.820 4.300 ;
        RECT 729.980 3.500 733.860 4.300 ;
        RECT 735.020 3.500 738.900 4.300 ;
        RECT 740.060 3.500 743.940 4.300 ;
        RECT 745.100 3.500 748.980 4.300 ;
        RECT 750.140 3.500 754.020 4.300 ;
        RECT 755.180 3.500 759.060 4.300 ;
        RECT 760.220 3.500 764.100 4.300 ;
        RECT 765.260 3.500 769.140 4.300 ;
        RECT 770.300 3.500 774.180 4.300 ;
        RECT 775.340 3.500 779.220 4.300 ;
        RECT 780.380 3.500 784.260 4.300 ;
        RECT 785.420 3.500 789.300 4.300 ;
        RECT 790.460 3.500 794.340 4.300 ;
        RECT 795.500 3.500 799.380 4.300 ;
        RECT 800.540 3.500 804.420 4.300 ;
        RECT 805.580 3.500 809.460 4.300 ;
        RECT 810.620 3.500 814.500 4.300 ;
        RECT 815.660 3.500 819.540 4.300 ;
        RECT 820.700 3.500 824.580 4.300 ;
        RECT 825.740 3.500 829.620 4.300 ;
        RECT 830.780 3.500 834.660 4.300 ;
        RECT 835.820 3.500 839.700 4.300 ;
        RECT 840.860 3.500 844.740 4.300 ;
        RECT 845.900 3.500 849.780 4.300 ;
        RECT 850.940 3.500 854.820 4.300 ;
        RECT 855.980 3.500 859.860 4.300 ;
        RECT 861.020 3.500 864.900 4.300 ;
        RECT 866.060 3.500 869.940 4.300 ;
        RECT 871.100 3.500 893.060 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 4.060 893.110 586.180 ;
      LAYER Metal4 ;
        RECT 117.740 21.930 175.540 288.870 ;
        RECT 177.740 21.930 252.340 288.870 ;
        RECT 254.540 21.930 329.140 288.870 ;
        RECT 331.340 21.930 405.940 288.870 ;
        RECT 408.140 21.930 482.740 288.870 ;
        RECT 484.940 21.930 559.540 288.870 ;
        RECT 561.740 21.930 629.860 288.870 ;
  END
END DSP48
END LIBRARY

