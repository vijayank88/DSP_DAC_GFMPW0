* NGSPICE file created from DSP48.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

.subckt DSP48 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] user_clock2 vdd vss wb_ACK wb_ADR[0] wb_ADR[10]
+ wb_ADR[11] wb_ADR[12] wb_ADR[13] wb_ADR[14] wb_ADR[15] wb_ADR[16] wb_ADR[17] wb_ADR[18]
+ wb_ADR[19] wb_ADR[1] wb_ADR[20] wb_ADR[21] wb_ADR[22] wb_ADR[23] wb_ADR[24] wb_ADR[25]
+ wb_ADR[26] wb_ADR[27] wb_ADR[28] wb_ADR[29] wb_ADR[2] wb_ADR[30] wb_ADR[31] wb_ADR[3]
+ wb_ADR[4] wb_ADR[5] wb_ADR[6] wb_ADR[7] wb_ADR[8] wb_ADR[9] wb_CYC wb_DAT_MISO[0]
+ wb_DAT_MISO[10] wb_DAT_MISO[11] wb_DAT_MISO[12] wb_DAT_MISO[13] wb_DAT_MISO[14]
+ wb_DAT_MISO[15] wb_DAT_MISO[16] wb_DAT_MISO[17] wb_DAT_MISO[18] wb_DAT_MISO[19]
+ wb_DAT_MISO[1] wb_DAT_MISO[20] wb_DAT_MISO[21] wb_DAT_MISO[22] wb_DAT_MISO[23] wb_DAT_MISO[24]
+ wb_DAT_MISO[25] wb_DAT_MISO[26] wb_DAT_MISO[27] wb_DAT_MISO[28] wb_DAT_MISO[29]
+ wb_DAT_MISO[2] wb_DAT_MISO[30] wb_DAT_MISO[31] wb_DAT_MISO[3] wb_DAT_MISO[4] wb_DAT_MISO[5]
+ wb_DAT_MISO[6] wb_DAT_MISO[7] wb_DAT_MISO[8] wb_DAT_MISO[9] wb_DAT_MOSI[0] wb_DAT_MOSI[10]
+ wb_DAT_MOSI[11] wb_DAT_MOSI[12] wb_DAT_MOSI[13] wb_DAT_MOSI[14] wb_DAT_MOSI[15]
+ wb_DAT_MOSI[16] wb_DAT_MOSI[17] wb_DAT_MOSI[18] wb_DAT_MOSI[19] wb_DAT_MOSI[1] wb_DAT_MOSI[20]
+ wb_DAT_MOSI[21] wb_DAT_MOSI[22] wb_DAT_MOSI[23] wb_DAT_MOSI[24] wb_DAT_MOSI[25]
+ wb_DAT_MOSI[26] wb_DAT_MOSI[27] wb_DAT_MOSI[28] wb_DAT_MOSI[29] wb_DAT_MOSI[2] wb_DAT_MOSI[30]
+ wb_DAT_MOSI[31] wb_DAT_MOSI[3] wb_DAT_MOSI[4] wb_DAT_MOSI[5] wb_DAT_MOSI[6] wb_DAT_MOSI[7]
+ wb_DAT_MOSI[8] wb_DAT_MOSI[9] wb_SEL wb_STB wb_WE wb_clk_i wb_rst_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6209__A2 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3691__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5968__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3428__C1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _0068_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input108_I wb_DAT_MOSI[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6845_ _0153_ net65 dacArea_dac_cnt_3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6393__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6776_ dspArea_regP\[40\] _2942_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3988_ _0203_ net121 _0170_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _0219_ _3057_ _1811_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_17_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5658_ _0529_ _3101_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input73_I wb_ADR[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ _0799_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5589_ _0791_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4459__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5959__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A3 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3993__I0 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6136__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3673__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__B2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3869__I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4960_ _1039_ _1042_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4622__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ net105 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _1080_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6630_ _0792_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6375__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3842_ _3292_ _3331_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_34_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ _2723_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3773_ dacArea_dac_cnt_5\[5\] net40 _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4925__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5512_ _1695_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6127__A1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _2663_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6678__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5443_ _0180_ _3079_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5374_ _1456_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4325_ _0181_ _3029_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _0453_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5102__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4456__A4 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4187_ _0369_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6921__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6828_ _0136_ net65 dacArea_dac_cnt_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _2911_ _2913_ _2926_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_12_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3910__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4907__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4110_ _0285_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5090_ _0240_ _3017_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4041_ net98 net159 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_65_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _2076_ _0297_ _2172_ _1461_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_18_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _1131_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4071__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6348__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4874_ _1062_ _1063_ _1064_ _1057_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _2776_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3825_ dacArea_dac_cnt_7\[1\] net53 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_21_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5020__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ _2712_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ dacArea_dac_cnt_5\[1\] net36 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5571__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _2647_ _2648_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3687_ _3207_ _3209_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _1591_ _1593_ _1610_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5323__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5357_ _1440_ _1441_ _1439_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0207_ _3008_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ _1472_ _1473_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA_input36_I la_data_in[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7027_ net147 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ _0438_ _0392_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A1 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6817__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3948__I0 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6967__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5078__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5617__A3 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3610_ dacArea_dac_cnt_1\[2\] net2 _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_31_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5553__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _0713_ _0692_ _0783_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5583__B _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ dspArea_regA\[23\] _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3882__I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _0232_ _3075_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3472_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5211_ _1397_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6191_ _2317_ _2318_ _2316_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3867__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ dspArea_regP\[17\] _1228_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5069__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _3173_ _1162_ _1262_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4816__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4024_ _0233_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A3 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _2154_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_52_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4044__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5241__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4926_ _0364_ _3044_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5792__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _0876_ _0954_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3993__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ dacArea_dac_cnt_6\[4\] net48 _3302_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6741__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5544__A2 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3555__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _2649_ _2700_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3792__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3739_ dacArea_dac_cnt_4\[5\] net31 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _2334_ _2413_ _2486_ _2565_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5409_ _1508_ _1594_ _1517_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_79_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6389_ _2563_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A3 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5578__B _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _1844_ _1846_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5774__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _0900_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _1786_ _1794_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4642_ _0195_ _3032_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5526__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _0667_ _0669_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2348_ _2487_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3524_ dspArea_regP\[19\] _3004_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6243_ _0792_ _2419_ _2420_ _1461_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3455_ _3031_ net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ dspArea_regP\[28\] _2223_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5125_ _0406_ _3056_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _1242_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_73_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4007_ _0219_ net100 _0169_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5214__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _0177_ _3105_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4909_ _0206_ _3036_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5889_ _1960_ _1963_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5517__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3528__A1 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3700__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5453__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3464__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3464__C2 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5444__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6930_ _0084_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6861_ _0015_ net65 dacArea_dac_cnt_5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5812_ _1992_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6792_ _2949_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5743_ _1922_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5674_ _1741_ _1742_ _1739_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _0817_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4183__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _0200_ _3025_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3507_ _3071_ _3073_ net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3930__A1 _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4487_ _0592_ _0606_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _0241_ _3062_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3438_ dspArea_regP\[35\] _2992_ _3006_ _3017_ _3004_ dspArea_regP\[3\] _3018_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _2157_ _2160_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _1295_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _2182_ _2195_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5435__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5039_ dspArea_regP\[17\] _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4789__A3 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5738__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3980__I _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5674__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput120 wb_DAT_MOSI[6] net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5426__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4401__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4165__A1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _0592_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _1476_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _0470_ _0537_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _0173_ _3033_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6011_ _2187_ _2188_ _2189_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4468__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5417__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3428__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3428__C2 dspArea_regP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6090__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _0067_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _0152_ net65 dacArea_dac_cnt_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6775_ _2910_ _2859_ _2510_ _2941_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3987_ _0202_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _0213_ _3065_ _1696_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5657_ _0172_ _3097_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_15_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _0800_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5588_ dspArea_regP\[23\] _0259_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input66_I wb_ADR[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3903__A1 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4896__I _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ _0206_ _3019_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_46_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4459__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _2383_ _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5408__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3975__I _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__A1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6136__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__I1 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3910_ _3380_ _3371_ _3381_ _3373_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4890_ _1077_ _1078_ _1079_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ dacArea_dac_cnt_7\[4\] net57 _3330_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3885__I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3772_ _3275_ _3276_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6560_ _2725_ _2732_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5511_ _0205_ _3060_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6491_ _2581_ _2664_ _2663_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_8_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5442_ _0187_ _3075_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4689__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5373_ _1366_ _1453_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4324_ _0188_ _3025_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ _0203_ _3000_ _0408_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ _0383_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_28_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input120_I wb_DAT_MOSI[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _0135_ net65 dacArea_dac_cnt_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ _2924_ _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_7_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ _1879_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6689_ _0238_ _3102_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4129__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output172_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5629__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4301__A1 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4067__S _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6896__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__A1 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ _0246_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5991_ _2170_ _2171_ _0248_ _0790_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ dspArea_regP\[16\] _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6348__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _0786_ _0872_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ _2782_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3824_ _3142_ _3316_ _3317_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5020__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6543_ _2714_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3755_ _3173_ _3262_ _3263_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_20_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6474_ _2619_ _2623_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3686_ dacArea_dac_cnt_3\[2\] net19 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _1591_ _1593_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5323__A3 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5356_ _1440_ _1441_ _1439_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _0503_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _0236_ _3030_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7026_ net146 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4238_ _0324_ _0351_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input29_I la_data_in[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _0187_ _3012_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3948__I1 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3573__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__A1 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A3 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5078__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6027__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3540_ _3099_ _3100_ net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3564__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4761__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6911__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3471_ dspArea_regA\[10\] _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0205_ _3048_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6190_ _2317_ _2318_ _2316_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _1327_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5069__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5072_ _0792_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4023_ _0232_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5974_ _1998_ _2064_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4044__A3 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _0404_ _3041_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ _0965_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3807_ dacArea_dac_cnt_6\[4\] net48 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6741__A2 _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4787_ _0977_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _2696_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3555__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3738_ dacArea_dac_cnt_4\[5\] net31 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6457_ _1964_ _2070_ _2161_ _2260_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3669_ _3177_ _3196_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5408_ _1509_ _1510_ _1515_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6388_ _2506_ _2507_ _2562_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_47_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _0529_ dspArea_regA\[20\] _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6257__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4807__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A1 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _0901_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ _3173_ _1772_ _1873_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _0200_ _3029_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__A3 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4734__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ dspArea_regP\[11\] _0668_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6311_ _2351_ _2483_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3523_ _3086_ _2999_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3454_ dspArea_regP\[38\] _2992_ _3006_ _3030_ _3022_ dspArea_regP\[6\] _3031_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6242_ dspArea_regP\[29\] _0874_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _2349_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5613__I _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ _0364_ _3052_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5055_ _1110_ _1243_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ _0218_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6957__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _0186_ _3097_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _0210_ _3032_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5888_ _1980_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input96_I wb_ADR[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__I0 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4839_ _0935_ _0937_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5517__A3 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3528__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6190__A3 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _0972_ _3086_ _2580_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5150__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6650__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3464__A1 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3464__B2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5205__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6641__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5444__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3888__I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6860_ _0014_ net65 dacArea_dac_cnt_5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5811_ _1989_ _1990_ _1991_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6791_ _2951_ _2948_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5742_ _1923_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_31_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4007__I0 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _1820_ _1853_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__4707__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4624_ _0205_ _3024_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5380__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _0663_ _0747_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3506_ dspArea_regP\[16\] _3072_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3930__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _0602_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6225_ _2401_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5132__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3437_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _2176_ _2259_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5107_ _0206_ _3044_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ _2185_ _2194_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5435__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _0529_ _3074_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I la_data_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5738__A3 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5123__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3685__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput110 wb_DAT_MOSI[1] net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput121 wb_DAT_MOSI[7] net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A2 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A3 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4165__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _0474_ _0476_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4271_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ _2187_ _2188_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5665__A2 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input3_I la_data_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5417__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3428__A1 dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3428__B2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _0066_ clknet_3_1__leaf_wb_clk_i dspArea_regB\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6090__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6843_ _0151_ net65 dacArea_dac_cnt_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6774_ _0244_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5725_ _1904_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _1839_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _0724_ _0742_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5587_ _0355_ _1771_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3903__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4538_ _0210_ _3015_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input59_I la_data_in[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5105__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4469_ _0662_ _0663_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6208_ _2314_ _2384_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _0219_ _3076_ _2210_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_58_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6605__A1 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6081__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__A1 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3991__I _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5647__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _3328_ _3326_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_32_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5583__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ dacArea_dac_cnt_5\[4\] net39 _3273_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5510_ _0209_ _3056_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _2588_ _2589_ _2586_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5335__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5441_ _1616_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ _1360_ _1357_ _1454_ _1354_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _0512_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4254_ _0361_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3649__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4310__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ _0336_ _0384_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_27_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6063__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4074__A1 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input113_I wb_DAT_MOSI[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3821__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _0134_ net65 dacArea_dac_cnt_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _2921_ _2923_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5574__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3969_ _0187_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_17_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _1882_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6688_ _2855_ _2857_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _1821_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5629__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__I _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5565__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__I _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4766__B _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6840__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2167_ _2169_ _2161_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _0529_ _3068_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _0708_ _0709_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_36_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ _0243_ _3090_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3823_ dacArea_dac_cnt_7\[0\] net52 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6542_ _2656_ _2661_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3754_ _3260_ _3261_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5308__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6473_ _2614_ _2618_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3685_ _3177_ _3208_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5859__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _1595_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_12_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _1505_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6808__A1 dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4306_ _0455_ _0463_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5286_ _0972_ _3030_ _1394_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7025_ net145 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4237_ _0399_ _0433_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__4295__A1 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4168_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4047__A1 dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4099_ _0190_ _3001_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6809_ dspArea_regP\[45\] dspArea_regP\[44\] _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4770__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3494__C1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6027__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4589__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6092__I _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3470_ _3043_ net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5140_ dspArea_regP\[18\] _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6266__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _1252_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4816__A3 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5777__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ _2060_ _2063_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_18_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4924_ _0189_ _3050_ _1021_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5529__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _0966_ _1043_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3806_ _3292_ _3303_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4201__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4786_ _0241_ _3001_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6525_ _2697_ _2698_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3737_ _3234_ _3249_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _2629_ _2630_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3668_ dacArea_dac_cnt_2\[6\] net15 _3195_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5407_ _1492_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4504__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _2506_ _2507_ _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3599_ _3112_ _3141_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6886__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5338_ _0172_ _3085_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input41_I la_data_in[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6257__A2 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4268__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _1456_ _1361_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A3 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5940__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A1 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6420__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _0759_ _0831_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4734__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _0763_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6310_ _2351_ _2483_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3522_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6241_ _2413_ _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3453_ _3029_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6172_ _2271_ _2283_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5123_ _0404_ _3049_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5054_ _1143_ _1144_ _1142_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _0217_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ dspArea_regP\[26\] _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _0217_ _3029_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_16_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5887_ _1983_ _2065_ _2068_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__4973__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _1023_ _1027_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4025__I1 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input89_I wb_ADR[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A1 dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0299_ _0960_ _0961_ _0157_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6508_ _0229_ _3094_ _2521_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_20_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _2597_ _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3449__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3464__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6901__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6402__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6641__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5810_ _1989_ _1990_ _1991_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6790_ _2944_ _2950_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__4404__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5741_ _0406_ _3084_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4955__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ _1854_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4007__I1 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4623_ _0209_ _3019_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_15_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5904__A1 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3409__I _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4554_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3505_ _3003_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4485_ _0604_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6224_ _0237_ _3066_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3436_ _3015_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5132__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _2268_ _2331_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _0210_ _3040_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _2173_ _0297_ _2265_ _1461_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6924__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5037_ _0173_ _3069_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4643__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6396__A1 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _2118_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4946__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5123__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5674__A3 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput100 wb_DAT_MOSI[10] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput111 wb_DAT_MOSI[20] net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput122 wb_DAT_MOSI[8] net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4634__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5362__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4270_ _0465_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6947__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3899__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3428__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _0065_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6090__A3 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6842_ _0150_ net65 dacArea_dac_cnt_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6773_ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4928__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3985_ _0200_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ _1905_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _1835_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4606_ _0728_ _0741_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_50_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ dspArea_regP\[22\] _1770_ _0441_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4537_ _0217_ _3012_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5105__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _0178_ _3041_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6207_ _2209_ _2380_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3419_ _3001_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4399_ _0174_ _3041_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3667__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6138_ _0213_ _3086_ _2110_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6605__A2 _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _2245_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__A1 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A3 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ dacArea_dac_cnt_5\[4\] net39 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6780__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__A2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3594__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ _1624_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6532__A1 dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5335__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _1556_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4322_ _0515_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5099__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4253_ _0364_ _3011_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_45_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5902__I _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4184_ _0340_ _0342_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4310__A3 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input106_I wb_DAT_MOSI[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _0133_ net65 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6756_ _2921_ _2923_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3968_ _0186_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_17_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ _1888_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6687_ dspArea_regP\[37\] _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3899_ net101 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5638_ _0203_ _3066_ _1715_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5326__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input71_I wb_ADR[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _1752_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A3 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5262__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__I _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _0172_ _3065_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _0555_ _0559_ _0618_ _0694_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5005__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _2780_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3822_ dacArea_dac_cnt_7\[0\] net52 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _2652_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3753_ _3260_ _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6505__A1 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _2631_ _2642_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5308__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3684_ dacArea_dac_cnt_3\[2\] net19 _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _1600_ _1605_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ _1537_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ _0502_ _0462_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _0229_ _3038_ _1291_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4819__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7024_ net144 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4236_ _0357_ _0434_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5492__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _0360_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4098_ _0283_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4047__A2 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6808_ dspArea_regP\[45\] _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _2904_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3494__B1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3494__C2 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3997__I _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5538__A2 dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3549__A1 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5070_ _1254_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_1_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4021_ dspArea_regB\[13\] _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_49_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5226__A1 _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _2096_ _2149_ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _0183_ _3058_ _0928_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5529__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ _0887_ _1044_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ dacArea_dac_cnt_6\[4\] net48 _3302_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_4785_ _0975_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4201__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3736_ dacArea_dac_cnt_4\[5\] net31 _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6524_ _2601_ _2612_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3667_ dacArea_dac_cnt_2\[5\] net14 _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6455_ _2624_ _2628_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5406_ _1497_ _1500_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6386_ _2555_ _2558_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3598_ net143 net62 _3140_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__5701__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5337_ _1520_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5268_ _1350_ _1353_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input34_I la_data_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4268__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ _0167_ _3033_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _1298_ _1301_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5940__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6830__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A2 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ dspArea_regP\[12\] _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A2 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3942__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _3084_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _2414_ _2344_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3452_ _3028_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4498__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6171_ _2274_ _2282_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _0189_ _3058_ _1224_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5447__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5053_ _1143_ _1144_ _1142_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ _0216_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_66_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ dspArea_regP\[25\] _0173_ _3105_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _1093_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5886_ _1892_ _2066_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _0932_ _0934_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_14_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ dspArea_regP\[14\] _0299_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5922__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6507_ _2678_ _2679_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3933__A1 _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3719_ dacArea_dac_cnt_4\[1\] net27 _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _0839_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _2601_ _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _2543_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5438__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3449__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3449__C2 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3515__I _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6876__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ _0364_ _3079_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6157__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _1720_ _1738_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ _0217_ _3016_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4553_ _0182_ _0178_ _3041_ _3037_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_7_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3504_ _3070_ _2999_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ _0526_ _0535_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6223_ _2204_ _2375_ _2400_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3435_ dspArea_regA\[3\] _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _2179_ _2258_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4340__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _0217_ _3037_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6085_ _0296_ _2263_ _2264_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6093__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6632__A3 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4643__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6396__A2 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6471__I dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _2098_ _2100_ _2117_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5869_ _1939_ _1941_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3906__A1 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput101 wb_DAT_MOSI[11] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 wb_DAT_MOSI[21] net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput123 wb_DAT_MOSI[9] net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6899__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6139__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4322__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5822__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6910_ _0064_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6841_ _0149_ net65 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4389__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6772_ _2937_ _2938_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3984_ dspArea_regB\[7\] _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5723_ _0206_ _3068_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5654_ _1836_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5889__A1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4605_ _0644_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5585_ _1759_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4536_ _0729_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4467_ _0187_ _3033_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6206_ _2313_ _2315_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4313__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4398_ _0582_ _0593_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _2313_ _2314_ _2315_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _2135_ _2246_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _1207_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6057__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__A3 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6914__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _1366_ _1453_ _1350_ _1353_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_5_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4321_ _0516_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4252_ _0449_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4183_ _0340_ _0342_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6824_ _0132_ net65 dacArea_dac_cnt_0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6755_ _2895_ _2898_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3967_ dspArea_regB\[4\] _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3585__A2 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _0240_ _3042_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4782__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _0234_ _3106_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ _3370_ _3371_ _3372_ _3373_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5637_ _0198_ _3076_ _1621_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4534__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _1589_ _1654_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input64_I la_data_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4519_ _0685_ _0688_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5499_ _1605_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6211__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6937__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6762__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4828__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6450__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _1049_ _1056_ _1057_ _1058_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6202__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3821_ _3112_ _3315_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6540_ _2655_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3752_ dacArea_dac_cnt_5\[1\] net36 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6471_ dspArea_regP\[33\] _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3683_ _3206_ _3205_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5422_ _1606_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4516__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _1422_ _1538_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4304_ _0458_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5284_ _1470_ _1404_ _1407_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4819__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ net143 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4235_ _0388_ _0391_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5492__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4166_ _0363_ _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4097_ _0178_ _3012_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4047__A3 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6807_ dspArea_regP\[44\] _0298_ _2958_ _2963_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_23_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4999_ _0231_ _3020_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6738_ _2878_ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_23_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _2787_ _2790_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output170_I net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3494__A1 dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__B2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5235__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3549__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__I0 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4020_ _0215_ _0230_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_46_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5226__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _2022_ _2150_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_53_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4985__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4922_ _1111_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__I0 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _0947_ _0950_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3804_ _3300_ _3298_ _3301_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4784_ _0971_ _0973_ _0974_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4201__A3 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _2604_ _2611_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3735_ _3246_ _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6454_ _2624_ _2628_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3666_ _3193_ _3191_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _1497_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _2559_ _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3597_ _3138_ _3136_ _3139_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5701__A3 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5336_ _1521_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5267_ _1350_ _1353_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _0174_ _3030_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5198_ _1298_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input27_I la_data_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4149_ _0347_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6414__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3703__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4019__I0 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3520_ dspArea_regA\[19\] _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3942__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ dspArea_regA\[6\] _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6170_ _2268_ _2331_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5121_ _0183_ _3065_ _1127_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5447__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _1206_ _1238_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_38_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4003_ dspArea_regB\[10\] _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_66_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__A3 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _2123_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _1094_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5885_ _1951_ _1954_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4836_ dspArea_regP\[14\] _0933_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4767_ _0955_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6506_ _2572_ _2591_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3718_ _3110_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3933__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _0889_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6437_ _2604_ _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3649_ _3177_ _3180_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6368_ _2435_ _2450_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5319_ _0198_ _3062_ _1314_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_29_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _2391_ _2394_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5438__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3449__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3449__B2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3621__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4120__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5429__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__I dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _1733_ _1737_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _0812_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5365__A1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4552_ _0662_ _0664_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_15_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3503_ _3069_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4483_ _0661_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6222_ _2308_ _2311_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3434_ _3014_ net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ _2254_ _2257_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4340__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _1289_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _2260_ _2262_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5035_ _1221_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3441__I _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6820__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5937_ _2098_ _2100_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__3603__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _1939_ _1941_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_16_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input94_I wb_ADR[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6970__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _0406_ _3044_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5799_ _1882_ _1890_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3906__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A2 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 wb_DAT_MOSI[12] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput113 wb_DAT_MOSI[22] net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput124 wb_STB net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__A1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3842__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A3 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6139__A3 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3526__I dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4086__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6843__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _0148_ net65 dacArea_dac_cnt_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2914_ _2920_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3983_ _0166_ _0199_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4092__I dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _0210_ _3064_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5338__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _0176_ dspArea_regA\[21\] _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5916__I _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5889__A2 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _0227_ _3007_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5584_ _1766_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_15_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ _0227_ _3000_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3436__I _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4466_ _0182_ _3037_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6205_ _2379_ _2382_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3417_ dspArea_regA\[0\] _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5510__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _0178_ _3037_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _0207_ _3089_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6067_ _2142_ _2143_ _2141_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_46_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _0203_ _3042_ _1119_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _0123_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5329__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4001__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6866__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4068__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _0509_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4251_ _0207_ _3001_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4182_ _0375_ _0378_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA_input1_I la_data_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6048__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4059__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3806__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _0131_ net65 dacArea_dac_cnt_0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _2884_ _2899_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ _0166_ _0185_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5705_ _1886_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ dspArea_regP\[36\] _2813_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4782__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _3109_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ _1818_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4534__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _1651_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6889__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4518_ _0689_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _1608_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input57_I la_data_in[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6287__A2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5381__I dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _0643_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4298__A1 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _2231_ _2244_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5798__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4222__A1 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5722__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5789__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4461__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6202__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3820_ net150 net51 _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5894__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3751_ _3142_ _3259_ _3260_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5961__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _3111_ _2644_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ dacArea_dac_cnt_3\[1\] net18 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5421_ _0634_ _3045_ _1496_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5713__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5352_ _1435_ _1438_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ _0449_ _0450_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5283_ _1318_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ net151 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ _0388_ _0391_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4165_ _0328_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4096_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input111_I wb_DAT_MOSI[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4452__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _3112_ _2968_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4998_ _1113_ _1187_ _1122_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_23_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _2844_ _2905_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3949_ _0166_ _0171_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5952__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _2787_ _2790_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_20_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5619_ _0231_ _3045_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6599_ _2728_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3479__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6904__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6196__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__I1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _2057_ _2058_ _2054_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _0202_ _3038_ _1012_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4985__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _0947_ _0950_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__I1 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3803_ dacArea_dac_cnt_6\[3\] net47 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4783_ _0971_ _0973_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__4737__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _2691_ _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3734_ dacArea_dac_cnt_4\[4\] net30 _3244_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _2625_ _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3665_ dacArea_dac_cnt_2\[5\] net14 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5404_ _1500_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6384_ _2459_ _2460_ _2473_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3596_ dacArea_dac_cnt_0\[6\] net61 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5335_ _0177_ _3079_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_47_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6111__A1 _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _1366_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6927__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4217_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _1301_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _0284_ _0348_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_18_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4079_ _0184_ _3008_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4425__A1 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6178__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6350__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6102__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4019__I1 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _3027_ net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5144__A2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5120_ _1307_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5051_ _1239_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4655__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4002_ _3110_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ _2132_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4904_ _0221_ _3024_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5884_ _1951_ _1954_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6243__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3630__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5907__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _1024_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4766_ _0712_ _0956_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5383__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6505_ _2572_ _2591_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3717_ _3173_ _3232_ _3233_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4697_ _0815_ _0824_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6436_ _2609_ _2610_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6332__A1 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3648_ dacArea_dac_cnt_2\[2\] net10 _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6367_ _2436_ _2449_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3579_ _3118_ _3125_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3697__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4894__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5318_ _1503_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6298_ _2391_ _2394_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6635__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__A3 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5249_ _1330_ _1332_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3902__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3449__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4646__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5992__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5677__A3 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4620_ _0798_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4551_ _0744_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3502_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4482_ _0673_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6221_ _2303_ _2397_ _2398_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3433_ dspArea_regP\[34\] _2992_ _3006_ _3013_ _3004_ dspArea_regP\[2\] _3014_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _2327_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _1290_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ _2260_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4628__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _1222_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3851__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _2102_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4800__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5867_ _1935_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6553__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _0196_ _3040_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _1876_ _1959_ _1979_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input87_I wb_ADR[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4749_ _0938_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6419_ _2508_ _2512_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput103 wb_DAT_MOSI[13] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput114 wb_DAT_MOSI[23] net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput125 wb_WE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5044__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3542__I _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4086__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6770_ _2916_ _2919_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6783__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3982_ _0198_ net120 _0170_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ _0217_ _3061_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6535__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _0181_ _3089_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5338__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _0716_ _0795_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_15_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5583_ _1558_ _1559_ _1563_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4534_ _0223_ _3008_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _0650_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3416_ _2998_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6204_ _2380_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5510__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4396_ _0187_ _3029_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _0634_ _3080_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3452__I _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _2142_ _2143_ _2141_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6066__A3 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5274__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _0198_ _3050_ _1011_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_22_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ _0122_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ _2009_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6899_ _0053_ clknet_3_6__leaf_wb_clk_i dspArea_regA\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3512__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__A1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5017__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3537__I _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3751__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _0447_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _0379_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6960__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6822_ _0130_ net65 dacArea_dac_cnt_0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5559__A2 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2914_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ _0184_ net117 _0170_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__I _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _1883_ _1884_ _1885_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6508__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6684_ _2834_ _2837_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3896_ _3046_ _3360_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_17_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5635_ _1798_ _1800_ _1817_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3447__I _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _1652_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4517_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5497_ _1669_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _0223_ _3001_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4298__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4379_ _0574_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _2296_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _2137_ _2140_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6747__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6211__A3 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6833__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3750_ dacArea_dac_cnt_5\[0\] net35 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A2 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6779__S _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3681_ _3173_ _3204_ _3205_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_51_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _0213_ _3053_ _1398_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _1435_ _1438_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4302_ _0499_ _0491_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5282_ _1309_ _1319_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5477__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7021_ net150 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4233_ _0400_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_4_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _0364_ _3007_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _2998_ _0249_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4452__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input104_I wb_DAT_MOSI[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6805_ dspArea_regP\[44\] _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _1114_ _1115_ _1120_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6856__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _2850_ _2879_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3948_ _0168_ net99 _0170_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _2834_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3879_ _3346_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_30_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5618_ _1709_ _1801_ _1718_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6598_ _2761_ _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5549_ _1632_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3905__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3479__B1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3479__C2 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3640__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4131__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7022__I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6879__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _0197_ _3046_ _0919_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_64_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _0981_ _1039_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_61_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3802_ dacArea_dac_cnt_6\[3\] net47 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4782_ _0236_ _3009_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _2693_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3733_ dacArea_dac_cnt_4\[4\] net30 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6452_ _2626_ _2561_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3664_ _3177_ _3192_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5403_ _1576_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6383_ _2465_ _2472_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3595_ dacArea_dac_cnt_0\[6\] net61 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4370__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5334_ _0182_ _3074_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6111__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ _1369_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4216_ _0412_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _1371_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4147_ _0312_ _0314_ _0311_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3460__I _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _0184_ _3002_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4425__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6178__A2 dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4189__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3936__A1 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _0243_ _3102_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6350__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6102__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5144__A3 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7017__I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4104__A1 dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1124_ _1141_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4001_ _0166_ _0214_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5852__A1 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4655__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _2125_ _2126_ _2131_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4903_ _0226_ _3019_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5883_ _1998_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4834_ dspArea_regP\[15\] _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5907__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4765_ _0871_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6504_ _2575_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3716_ _3230_ _3231_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4696_ _0820_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6435_ _0242_ _3076_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3455__I _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3647_ _3178_ _3176_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6366_ _2540_ _2541_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3578_ dacArea_dac_cnt_0\[3\] net34 _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_5317_ _1483_ _1485_ _1502_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _2461_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6096__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _1330_ _1332_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input32_I la_data_in[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _1272_ _1280_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3909__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6571__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4885__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6087__A1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5834__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3860__A3 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4550_ _0655_ _0658_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3501_ dspArea_regA\[16\] _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _0674_ _0675_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6220_ _2305_ _2306_ _2320_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4325__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_143_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6586__I dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _2196_ _2328_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _0221_ _3032_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _2261_ _2171_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0176_ _3064_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6250__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ _2107_ _2112_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4800__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5866_ _2041_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_55_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0201_ _3038_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6553__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _1955_ _1958_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5356__A3 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4564__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _0847_ _0939_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4679_ _0794_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4316__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _2571_ _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _0211_ _3097_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput104 wb_DAT_MOSI[14] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput115 wb_DAT_MOSI[24] net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput126 wb_rst_i net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5816__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5807__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7030__I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3981_ _0197_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _1899_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4794__A1 dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5651_ _0188_ _3085_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6535__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4602_ _0720_ _0782_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_30_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5582_ _1553_ _1554_ _1660_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_8_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _0726_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _0654_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6203_ _0207_ _3093_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3415_ _2996_ _2997_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4395_ _0581_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _0212_ _3085_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _2231_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ _1204_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _0121_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ _2014_ _2017_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6898_ _0052_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5849_ _2029_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3908__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4537__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3512__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4528__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4000__I0 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7025__I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4700__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ dspArea_regP\[6\] _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_67_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6821_ _0129_ net65 dacArea_dac_cnt_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__I0 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6752_ _2916_ _2919_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_17_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3964_ _0183_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5703_ _1883_ _1884_ _1885_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6683_ _2830_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6508__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3895_ _3346_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ _1798_ _1800_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ _1505_ _1541_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3742__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4516_ _0707_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5496_ _1672_ _1680_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4447_ _0639_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3463__I _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _0219_ _3001_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6774__I _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _2228_ _2229_ _2227_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ dspArea_regP\[26\] _2136_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6747__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3733__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6435__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5410__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3680_ _3202_ _3203_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4921__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ _1519_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4301_ _0399_ _0492_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_47_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7020_ net148 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _0428_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ _0195_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6804_ _0250_ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ _1097_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6735_ _2900_ _2903_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3947_ _0169_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3458__I _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6666_ _2835_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3878_ net119 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _1710_ _1711_ _1716_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5165__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _2758_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4912__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ _1726_ _1730_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA_input62_I la_data_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5479_ _1579_ _1587_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3479__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3479__B2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6417__A1 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5069__B _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3403__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6950__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4131__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6408__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _0911_ _1040_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3801_ _3292_ _3299_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5395__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ _0972_ _3009_ _0898_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6520_ _2597_ _2613_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3732_ _3234_ _3245_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6451_ _2555_ _2558_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ dacArea_dac_cnt_2\[5\] net14 _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _1579_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6382_ _2557_ _2505_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3594_ _3118_ _3137_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5333_ _0188_ _3069_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4370__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5264_ _1448_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4215_ _0413_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5195_ _1374_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_9_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4146_ _0312_ _0314_ _0311_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _0178_ _3009_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6823__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4979_ _1081_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6718_ _0238_ _3106_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3936__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__I _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6649_ _0223_ _3106_ _2763_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_50_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6629__A1 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6846__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ _0213_ net123 _0170_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5852__A2 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3863__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4593__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5951_ _2125_ _2126_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_52_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _0231_ _3016_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5882_ _2060_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _0529_ _3064_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__A3 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _0797_ _0785_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _2573_ _2574_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3715_ _3230_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__3394__A3 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _0823_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6434_ _2607_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3646_ dacArea_dac_cnt_2\[1\] net9 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6365_ _0243_ _3066_ _2470_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3577_ dacArea_dac_cnt_0\[2\] net23 _3123_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5316_ _1483_ _1485_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2465_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__B _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6096__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__I _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _1428_ _1432_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _1266_ _1364_ _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA_input25_I la_data_in[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _0190_ _3008_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3909__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4031__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6869__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4098__A1 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5257__B _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7028__I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3500_ _3067_ net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _0599_ _0601_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3431_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4325__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5522__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _2250_ _2253_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _0226_ _3028_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _2157_ _2160_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5032_ _0180_ _3060_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5053__A3 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5934_ _2113_ _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4261__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5865_ _2043_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_61_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _0190_ _3046_ _0929_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4013__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5796_ dspArea_regP\[25\] _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4564__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _0851_ _0853_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4678_ _0797_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6417_ _2572_ _2576_ _2591_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_31_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3629_ dacArea_dac_cnt_1\[5\] net5 _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4316__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6348_ _0634_ _3093_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _2367_ _2389_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput105 wb_DAT_MOSI[15] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput116 wb_DAT_MOSI[2] net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6017__I _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5504__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5807__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4156__B _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _0196_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4243__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5650_ _1823_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4601_ _0720_ _0782_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5581_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4532_ _0650_ _0660_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4463_ _0655_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6202_ _0211_ _3089_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3414_ net92 _2988_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _0585_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _2308_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _2235_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _1184_ _1186_ _1203_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6966_ _0120_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4234__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _2014_ _2097_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5982__A1 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ _0051_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _0192_ dspArea_regA\[20\] _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input92_I wb_ADR[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _1862_ _1863_ _1861_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output179_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4473__A1 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5017__A3 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3433__C1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6191__B _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A2 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4528__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4000__I1 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__A3 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _0128_ net65 dacArea_dac_cnt_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6751_ _2917_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5964__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _0182_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _0236_ _3046_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6682_ _2833_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3894_ net100 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _1802_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4519__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__S _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _1682_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4515_ _0708_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ _1678_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4446_ _0640_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6692__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4377_ _0566_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_86_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _2226_ _2285_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__A2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6047_ _2225_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5247__A3 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4207__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5955__A1 dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _0103_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6435__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__C _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5946__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4153__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7036__I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4300_ _0445_ _0495_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6123__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ _1379_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4231_ _0369_ _0429_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6674__A2 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4162_ _0361_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4093_ _2998_ _0249_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_23_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6803_ _2936_ _2955_ _2964_ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4995_ _1102_ _1105_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _2901_ _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3946_ _2994_ _2986_ _2990_ _3345_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_17_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6665_ _2774_ _2785_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3877_ _3357_ _3347_ _3358_ _3350_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _1693_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5165__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _2766_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5547_ _1633_ _1635_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4912__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _1567_ _0297_ _1663_ _1461_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_input55_I la_data_in[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _0560_ _0617_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3479__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5928__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6353__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4903__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6408__A2 dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3890__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3559__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ dacArea_dac_cnt_6\[3\] net47 _3298_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4780_ _0233_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6592__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5395__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3731_ dacArea_dac_cnt_4\[4\] net30 _3244_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ _3189_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6450_ _2555_ _2558_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6344__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5401_ _1585_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6381_ _2556_ _2457_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3593_ dacArea_dac_cnt_0\[6\] net61 _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__3953__I0 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5332_ _1508_ _1518_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _1282_ _1449_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__A1 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4214_ _0177_ _3024_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5194_ _1380_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4145_ _0330_ _0343_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_68_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _0277_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_3_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3633__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _0244_ _3009_ _1082_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6717_ dspArea_regP\[38\] _2885_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3929_ _3109_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_50_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _2766_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5138__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _2629_ _2630_ _2701_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4897__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4649__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__A2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5594__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4360__I0 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _2127_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3615__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _1006_ _1091_ _1015_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_80_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5881_ _1916_ _2061_ _2062_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4832_ _0173_ _3061_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _0786_ _0872_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _2674_ _2675_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3714_ dacArea_dac_cnt_4\[1\] net27 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4694_ _0880_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _0238_ _3081_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3645_ _3110_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3953__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6364_ _2539_ _2469_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3576_ _3120_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3551__A1 dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _1487_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6295_ _2470_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6096__A3 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5172__C _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _1327_ _1329_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5177_ _1347_ _1348_ _1346_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3854__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4128_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6940__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I la_data_in[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4059_ _0174_ _3009_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6556__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6308__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5047__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__A1 dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ dspArea_regA\[2\] _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5522__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3533__A1 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5100_ _0231_ _3025_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _2176_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6963__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _0186_ _3057_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3836__A2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6786__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5933_ _0217_ _3065_ _2013_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3948__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4261__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6538__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5864_ _1936_ _1938_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _0184_ _3054_ _0844_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5795_ _0355_ _1977_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5210__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4746_ _0851_ _0853_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4677_ _0868_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ _2581_ _2586_ _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3628_ _3163_ _3161_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5513__A2 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3524__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _2519_ _2522_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3482__I _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3559_ _3109_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6278_ _2453_ _2454_ _2366_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xinput106 wb_DAT_MOSI[16] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput117 wb_DAT_MOSI[3] net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ _1415_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_76_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4019__S _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4252__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5201__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6836__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5504__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5268__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3818__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _0785_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ _1762_ _1764_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _0654_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _0656_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3506__A1 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ _0218_ _3085_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3413_ _2982_ _2985_ _2995_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4393_ _0586_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _2309_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _2239_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _1184_ _1186_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_39_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _0119_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5431__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6859__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _2017_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6896_ _0050_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _0195_ _3084_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3477__I _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5734__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5778_ _1862_ _1863_ _1861_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_6_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input85_I wb_ADR[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _0915_ _0916_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4101__I _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4170__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__I _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3433__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A2 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3433__C2 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4528__A3 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5489__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__I _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4161__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4464__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5661__A1 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _2886_ _2894_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3962_ _0181_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_56_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5964__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5701_ _0233_ _3046_ _1806_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _2850_ _2844_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3893_ _3368_ _3347_ _3369_ _3350_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5632_ _1807_ _1812_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5716__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3727__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5563_ _1744_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4514_ _0623_ _0624_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5494_ _0241_ _3034_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4445_ _0219_ _3000_ _0574_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6141__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4152__A1 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4376_ _0207_ _3012_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _2289_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2173_ _2222_ _2224_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_86_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5652__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4207__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _0102_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5955__A2 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3966__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _0033_ net65 dacArea_dac_cnt_7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output191_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4391__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4143__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5643__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5946__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4006__I _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3709__A1 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4382__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ _0383_ _0386_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6674__A3 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4685__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _0198_ _3000_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ dspArea_regP\[4\] _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ dspArea_regP\[43\] dspArea_regP\[42\] _2949_ _2956_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _1102_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6733_ _2872_ _2876_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3945_ _0167_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_20_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6664_ _2776_ _2784_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3876_ _3021_ _3348_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5615_ _1698_ _1701_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6595_ _2587_ _2710_ _0219_ _3106_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5546_ dspArea_regP\[21\] _1634_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5477_ _0792_ _1661_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4428_ _0561_ _0622_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_input48_I la_data_in[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3490__I _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4359_ _0555_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5625__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _0206_ _3084_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3939__A1 _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6353__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4364__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5092__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6041__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _3242_ _3240_ _3243_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3661_ dacArea_dac_cnt_2\[4\] net13 _3187_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6344__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4355__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _0241_ _3030_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6380_ _2452_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3592_ dacArea_dac_cnt_0\[5\] net56 _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5331_ _1516_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3953__I1 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5262_ _1342_ _1345_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5855__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _0181_ _3019_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ _0241_ _3021_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4144_ _0304_ _0344_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ _0263_ _0264_ _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_37_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input102_I wb_DAT_MOSI[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6032__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _1165_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6716_ dspArea_regP\[37\] _2856_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4594__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3928_ _3090_ _3383_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6647_ _2767_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6335__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3485__I _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3859_ net98 net125 net159 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_30_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6578_ _2630_ _2750_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5529_ _0406_ _3074_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A3 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4360__I1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4812__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _1007_ _1008_ _1013_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5880_ _1948_ _1949_ _1947_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__A1 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6892__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _0876_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6501_ _2609_ _2610_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _3142_ _3229_ _3230_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_18_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4693_ _0884_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6432_ _2605_ _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ _3173_ _3175_ _3176_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6363_ _2468_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3575_ dacArea_dac_cnt_0\[2\] net23 _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ _1492_ _1497_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__3551__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _0241_ _3066_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5828__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5245_ dspArea_regP\[18\] _1328_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ _1347_ _1348_ _1346_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_56_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _0327_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_68_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6253__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4058_ dspArea_regP\[2\] _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_37_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6556__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4319__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3943__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5819__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6244__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3781__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4030__I0 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3533__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5030_ _1209_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5038__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ _0211_ _3075_ _1906_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_53_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6538__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _1004_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5794_ dspArea_regP\[24\] _1976_ _0441_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5210__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4745_ _0931_ _0935_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_31_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ _0869_ _0796_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6415_ _2588_ _2589_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3627_ dacArea_dac_cnt_1\[5\] net5 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3524__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6346_ _2520_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_1_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3558_ net126 _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6277_ _2353_ _2362_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3489_ dspArea_regP\[45\] _2991_ _2998_ _3058_ _3022_ dspArea_regP\[13\] _3059_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xinput107 wb_DAT_MOSI[17] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput118 wb_DAT_MOSI[4] net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5228_ _0192_ _3060_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input30_I la_data_in[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5159_ _1182_ _1246_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4960__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4012__I0 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4712__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6465__A1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5268__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6217__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _0659_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _0192_ _3028_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6200_ _2374_ _2377_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3506__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ _2993_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4703__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4392_ _0587_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _0222_ _3075_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2232_ _2240_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_85_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _1188_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6964_ _0118_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5431__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _2083_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6895_ _0049_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5846_ _0404_ _3080_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4242__I0 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5777_ _1876_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3745__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4942__A1 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _0917_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input78_I wb_ADR[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3493__I _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4659_ _0763_ _0765_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6329_ _2458_ _2474_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4170__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5670__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3433__A1 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3433__B2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6953__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3736__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6686__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4161__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5110__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5661__A2 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _0180_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _0228_ _3054_ _1691_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _2849_ _2842_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3892_ _3042_ _3360_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5631_ _1813_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4924__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _1613_ _1745_ _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_8_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4513_ _0693_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5493_ _1676_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4444_ _0506_ _0636_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4152__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4375_ _0570_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _2224_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _2222_ _2224_ _2173_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5101__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6826__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6947_ _0101_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3488__I _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5955__A3 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6878_ _0032_ net65 dacArea_dac_cnt_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _0210_ _3068_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4915__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5340__A1 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3951__I _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5643__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6691__I1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3709__A2 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4382__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4022__I _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3861__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6849__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__A2 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _0193_ _3008_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_4_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _0215_ _0294_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _2963_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5398__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4993_ _1105_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6732_ _2867_ _2871_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3944_ dspArea_regB\[0\] _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4070__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6663_ _2830_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3875_ net118 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _1698_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ _2762_ _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_30_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ _1727_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5570__A1 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3972__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _1554_ _1568_ _1660_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_144_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _0562_ _0563_ _0616_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5322__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4358_ _0498_ _0500_ _0554_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_63_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _0368_ _0387_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5625__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _0210_ _3079_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3636__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5389__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4061__A1 dspArea_regP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6909__D _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__A1 dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4017__I _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6041__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3660_ dacArea_dac_cnt_2\[4\] net13 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3591_ _3134_ _3132_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5330_ _1509_ _1510_ _1515_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_6_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6388__B _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5261_ _1342_ _1345_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5855__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4212_ _0188_ _3016_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5192_ _1378_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4143_ _0308_ _0310_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6804__A1 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4074_ dspArea_regP\[2\] _0262_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _1073_ _1085_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6715_ _2863_ _2883_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3927_ net111 _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5791__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _2781_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3858_ net99 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5543__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _2649_ _2700_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3789_ _3288_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5528_ _0364_ _3069_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input60_I la_data_in[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _1627_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3857__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output147_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6023__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4337__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6262__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4273__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ _1018_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4576__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _0877_ _0951_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _2673_ _2608_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3712_ dacArea_dac_cnt_4\[0\] net26 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _0238_ _3002_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3643_ _3172_ _3174_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6431_ _0234_ _3081_ _2522_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5525__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6362_ _2534_ _2537_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3574_ _3118_ _3121_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5313_ _1498_ _1499_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6293_ _2468_ _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5828__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5244_ _1429_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5175_ _0355_ _1363_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4126_ _0193_ _3000_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_28_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _0168_ _3013_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4264__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5764__A1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _1086_ _1146_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4319__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _2797_ _2800_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5819__A2 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_230 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6244__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4255__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5755__A1 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6180__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4030__I1 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6483__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _2108_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5796__I dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ dspArea_regP\[24\] _0168_ dspArea_regA\[24\] _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4549__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _0203_ _3034_ _0920_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_61_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _1965_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4744_ _0848_ _0850_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4675_ _0778_ _0781_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3626_ _3118_ _3162_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6414_ _0219_ _3094_ _2527_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3557_ dspArea_regP\[31\] _3072_ net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6345_ _0222_ _3089_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6276_ _2353_ _2362_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_9_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput108 wb_DAT_MOSI[18] net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5227_ _0195_ _3056_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput119 wb_DAT_MOSI[5] net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _1242_ _1245_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_5_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input23_I la_data_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4109_ _0277_ _0279_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4237__A1 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _1276_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_38_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5985__A1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4012__I1 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4712__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6465__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6882__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4779__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A1 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _0364_ _3024_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3411_ net91 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5900__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _0193_ _3025_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4703__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6130_ _0227_ _3069_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A2 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ _0193_ _3097_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5012_ _1193_ _1198_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4219__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _0117_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _2086_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6894_ _0048_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5845_ _0188_ _3090_ _1934_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5195__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5776_ _1955_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4242__I1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4727_ _0918_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ dspArea_regP\[12\] _0764_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 wb_ADR[31] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3609_ _3148_ _3147_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4589_ _0713_ _0692_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6328_ _2458_ _2474_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _2358_ _2361_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_76_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3433__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__B _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6686__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4449__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ dspArea_regB\[3\] _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_51_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3891_ net123 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _0218_ _3053_ _1697_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6374__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4924__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5561_ _1648_ _1649_ _1645_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _0703_ _0704_ _0705_ _0706_ _0617_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_5492_ _1673_ _1674_ _1675_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__A2 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4443_ _0635_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4688__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4374_ _0512_ _0520_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _2287_ _2290_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _2124_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5101__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3663__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input125_I wb_WE vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _0100_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6877_ _0031_ net65 dacArea_dac_cnt_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6365__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _0216_ _3065_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5168__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input90_I wb_ADR[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ _1935_ _1939_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4915__A2 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output177_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6920__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6356__A1 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__I0 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3893__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ dspArea_regP\[3\] _0293_ _0259_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5095__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6800_ dspArea_regP\[43\] dspArea_regP\[42\] _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_63_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5398__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _1169_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6731_ _2884_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_16_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _3110_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4070__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6662_ _2831_ _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ _3355_ _3347_ _3356_ _3350_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5613_ _1701_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _2763_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5544_ dspArea_regP\[22\] _1728_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5475_ _1554_ _1568_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _0562_ _0563_ _0616_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5322__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4357_ _0498_ _0500_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3884__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4288_ _0451_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5086__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6943__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _0216_ _3075_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4833__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _0083_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5010__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__I _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5001__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4033__I _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ dacArea_dac_cnt_0\[5\] net56 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3872__I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5260_ _1384_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6966__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _0366_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _1375_ _1376_ _1377_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4142_ _0308_ _0310_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5068__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _0274_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3618__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4815__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4975_ _1076_ _1084_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6714_ _2865_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6423__I _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ _3391_ _3371_ _0154_ _3373_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5791__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _2782_ _2783_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3857_ _3112_ _3343_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6576_ _2649_ _2700_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5543__A2 dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3788_ dacArea_dac_cnt_6\[1\] net44 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3554__A1 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _0404_ _3065_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _1639_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input53_I la_data_in[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4409_ _0602_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _0244_ _3026_ _1477_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_75_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4282__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3957__I _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6839__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4054__S _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__I _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__I0 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4788__I _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3848__A2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4273__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5470__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4028__I _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _0803_ _0867_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5773__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3711_ dacArea_dac_cnt_4\[0\] net26 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3784__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _0882_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6430_ _0229_ _3090_ _2439_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ _3172_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5525__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6361_ _2535_ _2536_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3573_ dacArea_dac_cnt_0\[2\] net23 _3120_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ _0219_ _3042_ _1399_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _0237_ _3070_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5289__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5243_ dspArea_regP\[19\] _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3839__A2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5174_ dspArea_regP\[18\] _1362_ _0441_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ _0325_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6789__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _0253_ _0257_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6581__C _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5478__B _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5213__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _1003_ _1147_ _1148_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3909_ _3062_ _3360_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4889_ _1077_ _1078_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6628_ _2798_ _2755_ _2799_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6713__A1 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6559_ _2730_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_10_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_220 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_231 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_19_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4255__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3518__A1 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5691__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5930_ _2109_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3454__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__C2 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5861_ _1978_ _2042_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_55_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _0198_ _3042_ _0837_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_21_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5792_ _1971_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ dspArea_regP\[13\] _0849_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4674_ _0803_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6413_ _2444_ _2587_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3625_ dacArea_dac_cnt_1\[5\] net5 _3161_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6171__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _0227_ _3085_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3556_ dspArea_regP\[30\] _3072_ net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6275_ _2432_ _2451_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_88_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3487_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput109 wb_DAT_MOSI[19] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5226_ _0200_ _3053_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5682__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5157_ _1282_ _1342_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_56_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4108_ _0304_ _0308_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5987__I _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5088_ _1273_ _1274_ _1275_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input16_I la_data_in[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _2985_ _2995_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5985__A2 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5737__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6162__A2 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3920__A1 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3970__I _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6465__A3 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__I _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A3 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4400__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3410_ net88 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4164__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _0196_ _3020_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5900__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _0200_ _3089_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I la_data_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5011_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4219__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _0116_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5913_ _2092_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6893_ _0047_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _0183_ _3097_ _1837_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1796_ _1956_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4726_ _0192_ _3040_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ _0848_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_11_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput80 wb_ADR[22] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3608_ dacArea_dac_cnt_1\[1\] net64 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput91 wb_ADR[3] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4588_ _0716_ _0720_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6327_ _2492_ _2495_ _2502_ _2501_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3539_ dspArea_regP\[22\] _3004_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _2433_ _2387_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _0209_ _3044_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_76_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6189_ _2363_ _2366_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5958__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4449__A2 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4036__I _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _3366_ _3347_ _3367_ _3350_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_43_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3875__I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _1648_ _1649_ _1645_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_8_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4511_ _0623_ _0693_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5491_ _1673_ _1674_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__4137__A1 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4442_ _0636_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4688__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4373_ _0569_ _0519_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _0193_ _3101_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5637__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _0187_ _3105_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input118_I wb_DAT_MOSI[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _0099_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _0030_ net65 dacArea_dac_cnt_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5827_ _2005_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6365__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1841_ _1843_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4915__A3 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input83_I wb_ADR[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _0205_ _3028_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5689_ _1773_ _1871_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5876__A1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__I1 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4119__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _1172_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_23_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6730_ _2895_ _2898_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_1_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3942_ _0164_ _3348_ _0165_ _0157_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6895__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _2770_ _2786_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3873_ _3017_ _3348_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5612_ _1783_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6592_ _0223_ _3105_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5543_ _0529_ dspArea_regA\[22\] _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3581__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _1571_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4425_ dspArea_regP\[11\] _0259_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4356_ _0549_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4287_ _0482_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6283__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _2203_ _2205_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_74_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6035__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6928_ _0082_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6859_ _0013_ net65 dacArea_dac_cnt_5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5010__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6775__B _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6274__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5001__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3563__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _0403_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _1375_ _1376_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ _0336_ _0340_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6265__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4072_ dspArea_regP\[3\] _0275_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_49_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ _1070_ _1154_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6713_ _3110_ _2848_ _2882_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3925_ _3086_ _3383_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _2810_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5379__I0 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3856_ net151 net60 _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6575_ _2744_ _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3787_ _3142_ _3287_ _3288_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6740__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3554__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _0189_ _3076_ _1631_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6910__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5457_ _1640_ _1641_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4408_ _0527_ _0603_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6595__B _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5388_ _1572_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input46_I la_data_in[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _0474_ _0476_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ dspArea_regB\[14\] _3058_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4593__I1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6495__A1 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5222__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ _3112_ _3228_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ _0234_ _3001_ _0814_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3641_ dacArea_dac_cnt_2\[1\] net9 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6933__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _2432_ _2451_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4733__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3572_ _3119_ _3117_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5311_ _0213_ _3050_ _1296_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6291_ _2466_ _2467_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ _0529_ _3084_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _1354_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4124_ _0190_ _3001_ _0301_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_57_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 la_data_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4055_ _0215_ _0260_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input100_I wb_DAT_MOSI[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _1036_ _1037_ _1035_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3775__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3908_ net104 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4972__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _0236_ _3013_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3839_ dacArea_dac_cnt_7\[3\] net55 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6627_ _2744_ _2747_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_14_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _0242_ _3086_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _0216_ _3053_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6489_ _2588_ _2589_ _2586_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_10_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6477__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_210 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_221 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_232 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_59_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6229__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__I _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3518__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4191__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A1 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__A2 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6640__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3454__B2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3878__I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _0172_ dspArea_regA\[24\] _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _1257_ _1258_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4742_ _0932_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _0863_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6412_ _0213_ _3102_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3624_ _3159_ _3160_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6343_ _0232_ _3080_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3555_ dspArea_regP\[29\] _3072_ net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6274_ _2435_ _2450_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3486_ dspArea_regA\[13\] _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _0187_ _3061_ _1324_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5131__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6829__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1206_ _1343_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ _0274_ _0276_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5087_ _1273_ _1274_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5434__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ _0215_ _0245_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_25_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5198__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _2161_ _2167_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5370__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3920__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5122__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 wb_DAT_MISO[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6465__A4 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__A3 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5425__A2 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5189__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3739__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4936__A1 dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6689__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6677__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _0218_ _3029_ _1101_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5416__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _0115_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _0240_ _3050_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6892_ _0046_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _2023_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _1857_ _1860_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4725_ _0364_ _3036_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4656_ dspArea_regP\[13\] _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_11_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput70 wb_ADR[13] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3607_ _3111_ _3146_ _3147_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
Xinput81 wb_ADR[23] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _0778_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xinput92 wb_ADR[4] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6326_ _2500_ _2485_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3538_ _3098_ _2999_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6257_ _2383_ _2386_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3469_ dspArea_regP\[41\] _2992_ _3006_ _3042_ _3022_ dspArea_regP\[9\] _3043_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A2 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _0216_ _3040_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6188_ _2364_ _2294_ _2365_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5139_ _0529_ _3079_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4091__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3981__I _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3914__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5894__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4385__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _0623_ _0693_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5490_ _0237_ _3038_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_7_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4441_ _0206_ _3015_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5334__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3891__I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5885__A2 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4372_ _0515_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3896__A1 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _0200_ _3093_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _2220_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5637__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _0098_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__B _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ _0029_ net65 dacArea_dac_cnt_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__A1 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ _2006_ _2007_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4376__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ dspArea_regP\[23\] _1842_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4708_ _0209_ _3024_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5688_ _1866_ _1870_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input76_I wb_ADR[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _2482_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_89_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5628__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3639__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4064__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3811__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5316__A1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6816__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6292__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6044__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _1178_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _3106_ _3383_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ _2761_ _2769_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3872_ net117 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5611_ _1786_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6591_ _0228_ _3102_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _0172_ _3093_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5307__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _1574_ _1655_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4424_ _0355_ _0620_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4355_ _0551_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__A1 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4286_ _0411_ _0483_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_58_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6283__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _2186_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4294__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _0081_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4597__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _0012_ net65 dacArea_dac_cnt_5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _0237_ _3050_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5546__A1 dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _0792_ _2953_ _2954_ _3109_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4140_ _0305_ _0307_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _0168_ _3017_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6862__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4276__A1 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3484__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4973_ _1150_ _1153_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6712_ _0259_ _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3924_ net109 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ dspArea_regP\[36\] _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5379__I1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3855_ _3340_ _3338_ _3341_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6574_ _2745_ _2746_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3786_ dacArea_dac_cnt_6\[0\] net43 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _0183_ _3085_ _1522_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5456_ _1528_ _1530_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4407_ _0532_ _0534_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5700__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _1468_ _1480_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6595__C _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _0527_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input39_I la_data_in[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4269_ _0466_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_41_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4267__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6008_ _0233_ _3058_ _2106_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_46_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5519__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6495__A2 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6885__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4258__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _3110_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ dacArea_dac_cnt_0\[1\] net12 _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4733__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _1493_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_6_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _0972_ _3070_ _2377_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6486__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5241_ _0172_ _3080_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5172_ _1066_ _1355_ _1357_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_9_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _0184_ _3013_ _0281_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3404__I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 la_data_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4054_ dspArea_regP\[1\] _0258_ _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5997__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _1036_ _1037_ _1035_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3907_ _3378_ _3371_ _3379_ _3373_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_32_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4972__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _0233_ _3013_ _0989_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6174__A1 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _2748_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3838_ dacArea_dac_cnt_7\[3\] net55 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _2728_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5921__A1 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _3234_ _3274_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _1689_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6488_ _2656_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6477__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _1617_ _1618_ _1623_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XDSP48_200 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_211 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_222 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_233 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output145_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5988__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3917__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5912__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4715__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5979__A1 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6640__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__I0 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6900__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4810_ _0982_ _0983_ _1000_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A1 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5790_ _1972_ _1561_ _1767_ _1966_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ dspArea_regP\[14\] _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3894__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6156__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _0743_ _0864_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _2584_ _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3623_ dacArea_dac_cnt_1\[4\] net4 _3157_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5903__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6342_ _2423_ _2424_ _2427_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3554_ dspArea_regP\[28\] _3072_ net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3485_ _3055_ net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6273_ _2436_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5224_ _0182_ _3069_ _1223_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _1239_ _1240_ _1238_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4106_ dspArea_regP\[3\] _0275_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5086_ _0236_ _3021_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6631__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4037_ _0244_ net105 _0169_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4642__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6395__A1 dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _1971_ _1974_ _2168_ _1965_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4939_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6609_ _2777_ _2778_ _2779_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5370__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4849__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 net180 wb_DAT_MISO[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput191 net191 wb_DAT_MISO[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6923__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3979__I _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4633__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5189__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6138__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6689__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5113__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6960_ _0114_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _2090_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6891_ _0045_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _0202_ _3076_ _1925_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_62_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5773_ _1857_ _1860_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4927__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__I _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4724_ _0404_ _3033_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4655_ _0167_ _3057_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 la_data_in[63] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3606_ _3144_ _3145_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput71 wb_ADR[14] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput82 wb_ADR[24] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _0647_ _0779_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput93 wb_ADR[5] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6325_ _2500_ _2485_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3537_ _3097_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6256_ _2378_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3468_ _3041_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6946__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5207_ _1391_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6187_ _2226_ _2285_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3399_ _2977_ _2981_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4863__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _0173_ _3075_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input21_I la_data_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _1257_ _1258_ _1159_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_26_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3930__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__I _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4909__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6819__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _0210_ _3011_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6531__A1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _0505_ _0565_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3896__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6110_ _2240_ _2286_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _0188_ _3101_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _0097_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6874_ _0028_ net65 dacArea_dac_cnt_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__A2 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5825_ _0221_ _3060_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5756_ _1936_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3584__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4707_ _0216_ _3019_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5687_ _1866_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_11_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5325__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _0182_ _0177_ _3045_ _3041_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA_input69_I wb_ADR[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4569_ _0167_ _3053_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3887__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _2351_ _2483_ _2484_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _2415_ _2416_ _2333_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_58_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4836__A1 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6589__A1 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4064__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6761__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3992__I _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6513__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5316__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4827__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ net115 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ _3353_ _3347_ _3354_ _3350_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_31_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5004__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _1792_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6590_ _0234_ _3098_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ _1481_ _1656_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4423_ dspArea_regP\[10\] _0619_ _0441_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4354_ _0493_ _0491_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6807__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4285_ _0424_ _0427_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4818__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _0221_ _3068_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5491__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input123_I wb_DAT_MOSI[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5243__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _0080_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6857_ _0011_ net65 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _0234_ _3050_ _1902_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_50_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6788_ dspArea_regP\[41\] _0874_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5546__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3557__A1 dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5739_ _0404_ _3075_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_13_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output175_I net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4809__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4285__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3987__I _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6363__I _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3548__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4070_ _0174_ _3013_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5473__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3484__B1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3484__C2 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5225__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ dspArea_regP\[17\] _0259_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_45_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5776__A2 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _2851_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3787__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3923_ _3389_ _3371_ _3390_ _3373_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_20_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _2811_ _2812_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ dacArea_dac_cnt_7\[6\] net59 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5528__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3539__A1 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _2696_ _2699_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3785_ dacArea_dac_cnt_6\[0\] net43 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ _1707_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _1528_ _1530_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4406_ _0532_ _0534_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5700__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ _1471_ _1479_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4337_ _0532_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_8_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4268_ _0176_ _3028_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _2007_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ _0347_ _0350_ _0392_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_55_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3600__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _0063_ clknet_3_7__leaf_wb_clk_i dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A2 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4258__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3510__I _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3570_ _3110_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_10_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3941__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__S _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5694__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4497__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5171_ _1164_ _1358_ _1359_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4122_ _0317_ _0316_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4053_ _0250_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_37_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 la_data_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5997__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _1110_ _1142_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3906_ _3058_ _3360_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4886_ _0227_ _3021_ _0897_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _2795_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3837_ _3292_ _3327_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6174__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _0237_ _3090_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3768_ dacArea_dac_cnt_5\[4\] net39 _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_69_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3932__A1 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _1690_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6487_ _2657_ _2660_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3699_ dacArea_dac_cnt_3\[5\] net22 _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ _1617_ _1618_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA_input51_I la_data_in[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_201 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_212 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_223 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ _1366_ _1453_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_234 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5988__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6852__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5912__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__A1 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3933__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3505__I _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5428__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _0167_ _3060_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ _0775_ _0776_ _0774_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6410_ _0219_ _3098_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3622_ dacArea_dac_cnt_1\[4\] net4 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6341_ _2514_ _2515_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3553_ dspArea_regP\[27\] _3072_ net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _2441_ _2446_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3484_ dspArea_regP\[44\] _2991_ _2998_ _3054_ _3022_ dspArea_regP\[12\] _3055_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5223_ _1409_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_9_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5154_ _1239_ _1240_ _1238_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4105_ _0305_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_69_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ _0233_ _3021_ _1192_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_2_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4036_ _0243_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_72_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4642__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6395__A2 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5987_ _2070_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4938_ _1125_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input99_I wb_DAT_MOSI[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4869_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4158__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ _2777_ _2778_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_20_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _2710_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput170 net170 wb_DAT_MISO[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput181 net181 wb_DAT_MISO[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6138__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A3 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5821__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6898__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _2087_ _2088_ _2089_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_81_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6890_ _0044_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5841_ _0197_ _3085_ _1828_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _1892_ _1951_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4723_ _0189_ _3041_ _0845_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6129__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4654_ _0173_ _3053_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput50 la_data_in[54] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3605_ _3144_ _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
Xinput61 la_data_in[6] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput72 wb_ADR[15] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4585_ _0682_ _0683_ _0679_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput83 wb_ADR[25] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6324_ _2482_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput94 wb_ADR[6] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3536_ dspArea_regA\[22\] _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_143_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _2429_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_27_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3467_ _3040_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6301__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5206_ _1392_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6186_ _2226_ _2285_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3398_ _2978_ _2979_ _2980_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5137_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _0707_ _0710_ _0956_ _1256_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_input14_I la_data_in[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _0229_ net102 _0169_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__A1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A2 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4090__I0 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3593__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6531__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _0450_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _0182_ _3105_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I la_data_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _0096_ clknet_3_6__leaf_wb_clk_i dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_81_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6873_ _0027_ net65 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5824_ _0226_ _3056_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5022__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5755_ dspArea_regP\[24\] _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4706_ _0896_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4781__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5686_ _1867_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6913__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4637_ _0758_ _0760_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6522__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _0173_ _3049_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3519_ _3082_ _3083_ net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_1_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _2408_ _2411_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4499_ _0626_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6238_ _2268_ _2331_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4836__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _2327_ _2330_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6589__A2 _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4434__I _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6789__C _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3575__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6513__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4524__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4827__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ _3013_ _3348_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6201__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6936__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3566__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5540_ _1721_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_30_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _1542_ _1545_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4422_ _0560_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4353_ _0550_ _0490_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6807__A3 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4284_ _0424_ _0427_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4818__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6023_ _0231_ _3061_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3423__I _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4682__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input116_I wb_DAT_MOSI[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5243__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _0079_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _0010_ net65 dacArea_dac_cnt_4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ _0229_ _3058_ _1805_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4054__I0 dspArea_regP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _2950_ _2952_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3999_ _0212_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3557__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5738_ _0189_ _3086_ _1838_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I wb_ADR[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _1834_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_output168_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4809__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6959__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3548__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3936__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5170__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3484__A1 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3484__B2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _0355_ _1161_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_63_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _2878_ _2879_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3922_ _3081_ _3383_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4984__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ dacArea_dac_cnt_7\[6\] net59 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6641_ _0234_ _3102_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3539__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _2691_ _2695_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3784_ _3112_ _3286_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5523_ _0202_ _3062_ _1622_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__3418__I _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5454_ _1524_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _0595_ _0599_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__5161__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _1465_ _1569_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5700__A3 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4336_ _0471_ _0473_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4267_ _0181_ _3024_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6006_ _0225_ _3064_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_39_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4198_ _0356_ _0395_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6908_ _0062_ clknet_3_0__leaf_wb_clk_i dspArea_regB\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4975__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6839_ _0147_ net65 dacArea_dac_cnt_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3998__I _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5391__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3941__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5694__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _1167_ _1351_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _0318_ _0316_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_64_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6643__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5446__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _0253_ _0257_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 la_data_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ _1143_ _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3905_ net103 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _1075_ _0999_ _1002_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4709__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _2759_ _2760_ _2794_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3836_ dacArea_dac_cnt_7\[3\] net55 _3326_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_20_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3767_ _3271_ _3269_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6555_ _2726_ _2727_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5506_ _0221_ _3048_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3932__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3698_ _3217_ _3218_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _2658_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5134__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _1619_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_10_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XDSP48_202 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__5685__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_213 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5368_ _1553_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XDSP48_224 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_235 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_input44_I la_data_in[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4319_ _0193_ _3020_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5299_ _1412_ _1413_ _1418_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7038_ net151 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4948__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5373__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5125__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5428__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3521__I _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ _0775_ _0776_ _0774_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _3118_ _3158_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6340_ _2446_ _2448_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3552_ dspArea_regP\[26\] _3072_ net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3914__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _2315_ _2447_ _2382_ _2379_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__5116__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3483_ _3053_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _0201_ _3049_ _1315_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_9_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _1306_ _1338_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_9_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4104_ dspArea_regP\[4\] _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5084_ _0228_ _3030_ _1095_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _0242_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_49_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3431__I _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6742__I dspArea_regP\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _2164_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _1126_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _0965_ _1055_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _0238_ _3094_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4158__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5355__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3819_ _3312_ _3310_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4799_ _0216_ _3024_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _0219_ _3106_ _2582_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_14_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ dspArea_regP\[32\] _2643_ _0874_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5658__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput160 net160 wb_DAT_MISO[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3669__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput171 net171 wb_DAT_MISO[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output150_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput182 net182 wb_DAT_MISO[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4330__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6607__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6386__A3 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3516__I _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3832__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _2020_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5771_ _1820_ _1952_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ _0183_ _3049_ _0760_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4653_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput40 la_data_in[45] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3604_ dacArea_dac_cnt_1\[1\] net64 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xinput51 la_data_in[55] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 la_data_in[7] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _0682_ _0683_ _0679_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xinput73 wb_ADR[16] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput84 wb_ADR[26] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ dspArea_regP\[31\] _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput95 wb_ADR[7] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3535_ _3095_ _3096_ net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3426__I _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _2353_ _2362_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3466_ dspArea_regA\[9\] _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5205_ _0221_ _3036_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6185_ _2353_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3397_ net87 net86 net90 net89 _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_5136_ _1321_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _1050_ _1255_ _1256_ _0958_ _1059_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_42_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6842__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4018_ _0228_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5576__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2057_ _2058_ _2054_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_52_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4303__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3939__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5319__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4790__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4542__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6865__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A1 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6941_ _0095_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _0026_ net65 dacArea_dac_cnt_6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _0231_ _3053_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5754_ _0167_ dspArea_regA\[24\] _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _0881_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4781__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ _1766_ _1768_ _1868_ _1867_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _0828_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4567_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6306_ _2408_ _2411_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3518_ dspArea_regP\[18\] _3072_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4498_ _0623_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6286__A2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _2268_ _2331_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3449_ dspArea_regP\[37\] _2992_ _3006_ _3026_ _3022_ dspArea_regP\[5\] _3027_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_44_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ _3111_ _2346_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _0202_ _3046_ _1215_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4049__A1 dspArea_regP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6099_ _2275_ _2276_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4450__I _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6888__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6277__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5281__I _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5788__A1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4460__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6201__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4212__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5470_ _1542_ _1545_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5712__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4515__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4352_ _0451_ _0486_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6268__A2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4283_ _0464_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_59_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6022_ _2123_ _2201_ _2133_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6924_ _0078_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input109_I wb_DAT_MOSI[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6855_ _0009_ net65 dacArea_dac_cnt_4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5806_ _1987_ _1912_ _1915_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6786_ _2936_ _2944_ _2951_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3998_ _0211_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5951__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5737_ _0183_ _3093_ _1723_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4754__A2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _1848_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_input74_I wb_ADR[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4619_ _0222_ _3012_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5599_ _1782_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5276__I _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3469__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__A3 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3484__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__A1 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6422__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ dspArea_regP\[16\] _1160_ _0441_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4433__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3921_ net108 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4984__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _0229_ _3106_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3852_ _3292_ _3339_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6571_ _2740_ _2743_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5933__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ net148 net42 _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_5522_ _0197_ _3070_ _1513_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5453_ _1632_ _1636_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_12_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _0528_ _0531_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5384_ _1547_ _1548_ _1546_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ dspArea_regP\[8\] _0472_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3434__I _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4266_ _0187_ _3020_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6005_ _2184_ _2116_ _2119_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_41_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6661__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _0355_ _0397_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__A2 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5216__A3 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4424__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _0061_ clknet_3_0__leaf_wb_clk_i dspArea_regB\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _0146_ net65 dacArea_dac_cnt_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6177__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6769_ _2804_ _2931_ _2932_ _2935_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6390__I _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4120_ _0295_ _0297_ _0322_ _0157_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6643__A2 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4051_ _0255_ _0256_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4654__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 la_data_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _1017_ _1034_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _3376_ _3371_ _3377_ _3373_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6159__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4884_ _0923_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6623_ _2759_ _2760_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_32_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3835_ dacArea_dac_cnt_7\[2\] net54 _3325_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5906__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4709__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3429__I _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _0234_ _3090_ _2660_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3766_ dacArea_dac_cnt_5\[3\] net38 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _0226_ _3044_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ _0223_ _3097_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3697_ dacArea_dac_cnt_3\[4\] net21 _3215_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _1620_ _1621_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5134__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_203 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_214 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ _1550_ _1552_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_225 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__3696__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4318_ _0201_ _3012_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_43_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5298_ _1395_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input37_I la_data_in[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ net150 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4196__S _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4249_ _0366_ _0410_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5373__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6322__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3620_ dacArea_dac_cnt_1\[4\] net4 _3157_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5364__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3551_ dspArea_regP\[25\] _3072_ net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _0213_ _3094_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3482_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _0196_ _3057_ _1214_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4875__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _1339_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4103_ _0168_ _3020_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5083_ _1271_ _1202_ _1205_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4627__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _0241_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_42_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3850__A2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5985_ _1960_ _1963_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ dspArea_regB\[2\] _3060_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3602__A2 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _0871_ _0957_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6606_ _0234_ _3094_ _2709_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3818_ dacArea_dac_cnt_6\[6\] net50 _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4158__A3 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5355__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4798_ _0986_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _2706_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3749_ dacArea_dac_cnt_5\[0\] net35 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_4_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5107__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _2631_ _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5419_ _1601_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xoutput150 net150 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput161 net161 wb_DAT_MISO[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6399_ _2528_ _2530_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput172 net172 wb_DAT_MISO[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput183 net183 wb_DAT_MISO[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_87_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output143_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__I _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3532__I _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ _1854_ _1855_ _1853_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6782__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _0912_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6534__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _0842_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3603_ _3142_ _3143_ _3144_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xinput30 la_data_in[36] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput41 la_data_in[46] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput52 la_data_in[56] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _0743_ _0774_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xinput63 la_data_in[8] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6322_ _3111_ _2498_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput74 wb_ADR[17] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput85 wb_ADR[27] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3534_ dspArea_regP\[21\] _3004_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput96 wb_ADR[8] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ dspArea_regP\[29\] _2352_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3465_ _3039_ net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5204_ _0225_ _3032_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6184_ _2358_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ net74 net73 net76 net75 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_5135_ _1322_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3442__I _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5066_ _0955_ _1048_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4017_ _0227_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _2120_ _2145_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4919_ _1108_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5899_ _2077_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__A2 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3511__A1 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3814__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3527__I _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6940_ _0094_ clknet_3_7__leaf_wb_clk_i dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3805__A2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _0025_ net65 dacArea_dac_cnt_6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _1919_ _2003_ _1928_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6755__A1 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3569__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5753_ _0173_ _3101_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _0222_ _3015_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3865__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _1755_ _1758_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _0751_ _0754_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3437__I _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _0758_ _0759_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__5730__A2 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _2478_ _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _3081_ _2999_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4497_ _0689_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6236_ _2334_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3448_ _3025_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6167_ dspArea_regP\[28\] _2345_ _0441_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _0197_ _3053_ _1118_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _0236_ _3062_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _1137_ _1140_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__A2 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3732__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A1 dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5788__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4212__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5960__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _0561_ _0564_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5712__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4351_ _0501_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4282_ _0477_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_3_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4279__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _2125_ _2126_ _2131_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_67_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _0077_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6854_ _0008_ net65 dacArea_dac_cnt_4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _1832_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _2940_ _2943_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3997_ _0210_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_50_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _1917_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _1726_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _0232_ _3000_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ _1677_ _1781_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input67_I wb_ADR[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _0198_ _3030_ _0588_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6219_ _2305_ _2306_ _2320_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4442__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6855__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3469__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3469__C2 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4130__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3920_ _3387_ _3371_ _3388_ _3373_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_45_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ dacArea_dac_cnt_7\[6\] net59 _3338_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _2741_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3782_ _3283_ _3281_ _3284_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5933__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _1704_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _1525_ _1527_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ dspArea_regP\[9\] _0530_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5383_ _1547_ _1548_ _1546_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4334_ _0528_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5449__A1 dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4265_ _0455_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_86_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6004_ _2034_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4196_ dspArea_regP\[6\] _0396_ _0259_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3450__I _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input121_I wb_DAT_MOSI[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6878__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6906_ _0060_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _0145_ net65 dacArea_dac_cnt_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _2905_ _2933_ _2934_ _2924_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5924__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__A1 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _1900_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6699_ _2815_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output173_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4179__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6340__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4103__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ _0174_ _3002_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6067__B _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5851__A1 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4654__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 la_data_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4406__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _1030_ _1033_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3903_ _3054_ _3360_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ _0914_ _0924_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6622_ _2787_ _2790_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3834_ _3322_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5906__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3917__A1 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _0229_ _3098_ _2579_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3765_ dacArea_dac_cnt_5\[3\] net38 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5504_ _0231_ _3041_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6484_ _0227_ _3093_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3696_ dacArea_dac_cnt_3\[4\] net21 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5435_ _0406_ _3068_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__I _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1550_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_204 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_215 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_226 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4317_ _0513_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5297_ _1400_ _1403_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7036_ net148 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4248_ _0446_ _0409_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ _0168_ _3029_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4333__A1 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5833__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _3107_ _3108_ net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4572__A1 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3481_ dspArea_regA\[12\] _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4324__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _1406_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4875__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5151_ _1220_ _1237_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5480__I _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4102_ _0174_ _3017_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5082_ _1122_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4096__I _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4033_ _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_2_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1876_ _1959_ _2069_ _1979_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5052__A2 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _0180_ _3056_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4866_ _0955_ _1048_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6605_ _2659_ _2763_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6916__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3817_ dacArea_dac_cnt_6\[6\] net50 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4797_ _0987_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4563__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3748_ _3112_ _3258_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6536_ _2707_ _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _2639_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3679_ _3202_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__4315__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput140 net140 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5418_ _1602_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xoutput151 net151 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6398_ _2523_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput162 net162 wb_DAT_MISO[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput173 net173 wb_DAT_MISO[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput184 net184 wb_DAT_MISO[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5349_ _1532_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_43_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4000__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5815__A1 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4618__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ net147 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5291__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7020__I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6939__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3596__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _0835_ _0838_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _0843_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6534__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput20 la_data_in[27] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3602_ dacArea_dac_cnt_1\[0\] net63 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput31 la_data_in[37] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4545__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _0775_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput42 la_data_in[47] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 la_data_in[57] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput64 la_data_in[9] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6321_ dspArea_regP\[30\] _2497_ _0874_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput75 wb_ADR[18] net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3533_ _3094_ _2999_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 wb_ADR[28] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput97 wb_ADR[9] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6252_ dspArea_regP\[30\] _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ dspArea_regP\[40\] _2992_ _3006_ _3038_ _3022_ dspArea_regP\[8\] _3039_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5203_ _0231_ _3029_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6183_ _2290_ _2359_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3395_ net79 net78 net81 net80 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5134_ _0176_ _3068_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ _1056_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6470__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4016_ _0226_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_26_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _2146_ _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5586__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4918_ _1088_ _1090_ _1107_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ _2078_ _1997_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_16_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input97_I wb_ADR[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ _0944_ _0945_ _0943_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _2692_ _2596_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6289__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3511__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5264__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3578__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4775__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5295__I _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5255__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _0024_ net65 dacArea_dac_cnt_6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ _1920_ _1921_ _1926_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5752_ _1931_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4703_ _0232_ _3008_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3718__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _1755_ _1758_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4634_ _0197_ _3034_ _0657_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_11_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ _0177_ _3045_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6304_ _2479_ _2480_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3881__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3516_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4496_ _0690_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6235_ _2348_ _2412_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3447_ _3024_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3453__I _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _2334_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _1304_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6097_ _0233_ _3062_ _2205_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _1220_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I la_data_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6434__A1 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5237__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4350_ _0545_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4920__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4281_ _0417_ _0478_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6673__A1 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6020_ _2107_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input4_I la_data_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5228__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6922_ _0076_ clknet_3_6__leaf_wb_clk_i dspArea_regB\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _0007_ net65 dacArea_dac_cnt_4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5804_ _1823_ _1833_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__4739__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6784_ _2948_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ _0209_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5400__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5735_ _0202_ _3070_ _1829_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3448__I _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5666_ _1730_ _1732_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5164__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4617_ _0809_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5597_ _0242_ _3034_ _1678_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_11_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _0724_ _0742_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _0599_ _0601_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _2279_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _2250_ _2253_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3911__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6719__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3402__A1 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6655__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3469__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3469__B2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4130__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6407__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ dacArea_dac_cnt_7\[5\] net58 _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3781_ dacArea_dac_cnt_5\[6\] net41 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5933__A3 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5520_ _1684_ _1686_ _1703_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_9_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5451_ dspArea_regP\[20\] _1526_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _0596_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5382_ _1555_ _1564_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ dspArea_regP\[9\] _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5449__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ _0458_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6003_ _2025_ _2035_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4195_ _0356_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_39_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3880__A1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input114_I wb_DAT_MOSI[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _0059_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6836_ _0144_ net65 dacArea_dac_cnt_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _2911_ _2925_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3979_ _0195_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3935__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5718_ _0222_ _3056_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ _2810_ _2814_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _1831_ _1832_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_40_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A2 dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4179__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5376__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__I0 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3926__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5128__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4103__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5300__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5851__A2 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput7 la_data_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6800__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _1124_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3902_ net102 _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4882_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6621_ _2791_ _2792_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5367__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3833_ dacArea_dac_cnt_7\[2\] net54 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6552_ _2724_ _2666_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3917__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3764_ _3234_ _3270_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5503_ _1616_ _1687_ _1625_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5119__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__I0 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6483_ _0972_ _3090_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4590__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _3177_ _3216_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5434_ _0364_ _3065_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5365_ _1369_ _1452_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XDSP48_205 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_216 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_227 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_4316_ _0189_ _3021_ _0468_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5296_ _1400_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6095__A2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ net147 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4247_ _0403_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6845__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5842__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _0174_ _3026_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _0127_ net65 dacArea_dac_cnt_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4333__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6086__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5597__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6631__B _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3546__I dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7018__I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ _3051_ net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4324__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6868__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _1233_ _1236_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4101_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5081_ _1113_ _1123_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6321__I0 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4032_ dspArea_regB\[15\] _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5824__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A3 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5588__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _1980_ _2162_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _0186_ _3053_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4260__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _0965_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_21_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _2775_ _2716_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _3292_ _3311_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _0221_ _3019_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6535_ _0223_ _3102_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3747_ net147 net33 _3257_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4563__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6466_ _1974_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3678_ dacArea_dac_cnt_3\[1\] net18 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4315__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _0206_ _3056_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xoutput130 net130 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput141 net141 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6397_ _2421_ _2422_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput152 net152 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput163 net163 wb_DAT_MISO[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput174 net174 wb_DAT_MISO[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5348_ _1428_ _1533_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xoutput185 net185 wb_DAT_MISO[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_input42_I la_data_in[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4079__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _0243_ _3021_ _1380_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7018_ net146 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5815__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5579__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__A3 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4251__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5503__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5806__A2 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _0177_ _3048_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3601_ dacArea_dac_cnt_1\[0\] net63 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput10 la_data_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput21 la_data_in[28] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4545__A2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput32 la_data_in[38] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _0661_ _0678_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput43 la_data_in[48] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 la_data_in[58] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6320_ _2486_ _2496_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xinput65 user_clock2 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_3532_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xinput76 wb_ADR[19] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput87 wb_ADR[29] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput98 wb_CYC net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6251_ _2425_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3463_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_143_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5202_ _1309_ _1389_ _1318_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4848__A3 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _2241_ _2355_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3394_ net83 net82 net85 net84 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _0180_ _3064_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5064_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _0225_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _2036_ _2053_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4917_ _1088_ _1090_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5981__A1 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5897_ _1985_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4848_ _0944_ _0945_ _0943_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4779_ _0228_ _3017_ _0813_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ _2593_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6289__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6449_ _2619_ _2623_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4472__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__C1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6906__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7031__I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ _1903_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5751_ _1932_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4702_ _0893_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5682_ _1776_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _0807_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _0186_ _3036_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6303_ _2396_ _2406_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3515_ _3079_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4495_ _0568_ _0615_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6234_ _2351_ _2408_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_143_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6140__A1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3446_ dspArea_regA\[5\] _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6165_ _2337_ _2340_ _2343_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5116_ _1284_ _1286_ _1303_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _0223_ _3070_ _2186_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5047_ _1233_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5949_ _2128_ _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5954__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5706__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6131__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4445__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6198__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3420__A2 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6370__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5173__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7026__I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4280_ _0421_ _0423_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6673__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6086__B _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4436__A1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _0075_ clknet_3_6__leaf_wb_clk_i dspArea_regB\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _0006_ net65 dacArea_dac_cnt_4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _1887_ _1984_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6783_ dspArea_regP\[41\] _2947_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__4739__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ dspArea_regB\[9\] _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _0197_ _3081_ _1714_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _1730_ _1732_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4616_ _0744_ _0745_ _0756_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _1777_ _1779_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4547_ _0728_ _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_2_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4478_ _0595_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6217_ _0244_ _3058_ _2280_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ _3010_ net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6148_ _2284_ _2322_ _2326_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _2179_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3402__A2 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6655__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3469__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A3 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3780_ dacArea_dac_cnt_5\[6\] net41 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6591__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _1633_ _1635_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6343__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4401_ dspArea_regP\[10\] _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5381_ dspArea_regP\[21\] _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4332_ _0529_ _3040_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4263_ _0459_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_68_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6002_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4194_ _0392_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_68_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _0058_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3887__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3632__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input107_I wb_DAT_MOSI[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6835_ _0143_ net65 dacArea_dac_cnt_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _2878_ _2930_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5385__A2 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ dspArea_regB\[6\] _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ _0226_ _3052_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6697_ _2858_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_13_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5648_ _1824_ _1825_ _1830_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input72_I wb_ADR[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__I0 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _1550_ _1552_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__3699__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3871__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5073__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4423__I1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4887__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5533__B _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 la_data_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6800__A2 dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4950_ _1137_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3901_ _3374_ _3371_ _3375_ _3373_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ _0976_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6620_ _2723_ _2733_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3832_ _3292_ _3323_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _2662_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3763_ dacArea_dac_cnt_5\[3\] net38 _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_20_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _1617_ _1618_ _1623_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6482_ _2652_ _2655_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5119__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__I1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3694_ dacArea_dac_cnt_3\[4\] net21 _3215_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_12_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5433_ _0404_ _3061_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5364_ _1448_ _1451_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XDSP48_206 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_217 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_4315_ _0184_ _3030_ _0414_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XDSP48_228 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _1403_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7034_ net146 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4246_ _0398_ _0443_ _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A3 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4177_ _0337_ _0339_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3853__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6818_ _0126_ net65 dacArea_dac_cnt_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ dspArea_regP\[38\] _2885_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6794__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5597__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6631__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3562__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7034__I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4100_ _0301_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5080_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6321__I1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ _0215_ _0239_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_42_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A2 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1983_ _2158_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_18_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1113_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_61_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4260__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _1047_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ dacArea_dac_cnt_6\[6\] net50 _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6603_ _2712_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4795_ _0225_ _3015_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ _0227_ _3098_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3746_ _3255_ _3253_ _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _1967_ _1970_ _2637_ _2638_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3677_ _3142_ _3201_ _3202_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5416_ _0210_ _3052_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput131 net131 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6396_ dspArea_regP\[32\] _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xoutput142 net142 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput153 net153 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3523__A1 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput164 net164 wb_DAT_MISO[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5347_ _1432_ _1434_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput175 net175 wb_DAT_MISO[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3472__I _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput186 net186 wb_DAT_MISO[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5278_ _1462_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4079__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6962__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I la_data_in[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7017_ net145 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4229_ _0383_ _0386_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6776__A1 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4251__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3817__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4427__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7029__I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3600_ _3109_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6835__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput11 la_data_in[19] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput22 la_data_in[29] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4580_ _0673_ _0677_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput33 la_data_in[39] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 la_data_in[49] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 la_data_in[59] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3531_ dspArea_regA\[21\] _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_7_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput66 wb_ADR[0] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput77 wb_ADR[1] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput88 wb_ADR[2] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput99 wb_DAT_MOSI[0] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6250_ _2354_ _2357_ _2426_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3462_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5201_ _1310_ _1311_ _1316_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6181_ _2287_ _2291_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3393_ _2976_ net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5132_ _0186_ _3061_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5063_ _1155_ _1158_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3808__A2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4014_ dspArea_regB\[12\] _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_42_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5965_ _2048_ _2052_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_80_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4916_ _1092_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5896_ _1988_ _1996_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3467__I _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _1003_ _1035_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_20_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4778_ _0968_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3729_ dacArea_dac_cnt_4\[3\] net29 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6517_ _2672_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5497__A1 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6379_ _2538_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__A1 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6858__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3983__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__B1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__C2 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5412__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5750_ _0176_ dspArea_regA\[22\] _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _0830_ _0840_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_30_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5681_ _1780_ _1861_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_31_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4632_ _0811_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ _0181_ _3040_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6302_ _2399_ _2405_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_7_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3514_ dspArea_regA\[18\] _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4494_ _0611_ _0614_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6233_ _2284_ _2409_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3445_ _3023_ net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6164_ _1971_ _1974_ _2341_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5115_ _1284_ _1286_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _2273_ _2215_ _2218_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_58_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1130_ _1234_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5403__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5948_ _0192_ dspArea_regA\[21\] _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_40_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5879_ _1948_ _1949_ _1947_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_21_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5706__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3717__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4390__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4142__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4693__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4445__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5945__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5881__A1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4684__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3570__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6920_ _0074_ clknet_3_7__leaf_wb_clk_i dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6851_ _0005_ net65 dacArea_dac_cnt_4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _0244_ _3042_ _1888_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6782_ dspArea_regP\[41\] _2947_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3994_ _0166_ _0208_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _1914_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _1840_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4615_ _0750_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5595_ _1778_ _1681_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4546_ _0731_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4477_ _0666_ _0670_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_143_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3428_ dspArea_regP\[33\] _2992_ _3006_ _3009_ _3004_ dspArea_regP\[1\] _3010_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6216_ _2392_ _2321_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _2324_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__3480__I _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _2254_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5624__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _1217_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5927__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3938__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5918__A2 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6343__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7037__I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _0167_ _3044_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5380_ _0355_ _1566_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ dspArea_regB\[0\] _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__A1 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4262_ _0452_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6001_ _2091_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5854__A1 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4193_ _0324_ _0351_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_39_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6903_ _0057_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6834_ _0142_ net65 dacArea_dac_cnt_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6919__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _2809_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3977_ _0166_ _0194_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5716_ _0232_ _3049_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6696_ _2863_ _2865_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3475__I _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5647_ _1824_ _1825_ _1830_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_5578_ _1465_ _1569_ _1570_ _1659_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_input65_I user_clock2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4529_ _0722_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5845__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4820__A2 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4970__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 la_data_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6261__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _3050_ _3360_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _0242_ _3002_ _0977_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3831_ dacArea_dac_cnt_7\[2\] net54 _3322_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6550_ _2721_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3762_ dacArea_dac_cnt_5\[2\] net37 _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _1600_ _1685_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3693_ _3213_ _3211_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6481_ _2653_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5432_ _0189_ _3070_ _1523_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _1465_ _1546_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_207 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _0510_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XDSP48_218 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5294_ _1468_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XDSP48_229 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7033_ net145 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4245_ _0437_ _0439_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4176_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3898__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6252__A1 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__A1 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6817_ _0125_ clknet_3_0__leaf_wb_clk_i _zz_1_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6891__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ dspArea_regP\[39\] _2915_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _2838_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4318__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4030__S _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5818__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6243__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6794__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4004__I _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _0238_ net104 _0169_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5285__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5037__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1983_ _2158_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_53_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4796__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ _1121_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4863_ _3173_ _0962_ _1054_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _2772_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4548__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ dacArea_dac_cnt_6\[5\] net49 _3309_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_32_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ dspArea_regB\[13\] _3011_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _0972_ _3094_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3745_ dacArea_dac_cnt_4\[6\] net32 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3771__A2 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6464_ _2634_ _2637_ _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3676_ dacArea_dac_cnt_3\[0\] net17 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5415_ _0217_ _3049_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6395_ dspArea_regP\[31\] _2511_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xoutput132 net132 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput143 net143 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput154 net154 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3523__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput165 net165 wb_DAT_MISO[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5346_ _1432_ _1434_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput176 net176 wb_DAT_MISO[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput187 net187 wb_DAT_MISO[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5277_ _1463_ _1383_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ net144 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4228_ _0411_ _0424_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input28_I la_data_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ _0358_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6225__A1 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4025__S _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6464__A1 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 la_data_in[1] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 la_data_in[2] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput34 la_data_in[3] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput45 la_data_in[4] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3530_ _3091_ _3092_ net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4950__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput56 la_data_in[5] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput67 wb_ADR[10] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput78 wb_ADR[20] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput89 wb_ADR[30] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3461_ dspArea_regA\[8\] _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5200_ _1293_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3392_ net124 _zz_1_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6180_ _2354_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5131_ _1309_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _1164_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _0215_ _0224_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5964_ _2135_ _2141_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _1097_ _1102_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_5895_ dspArea_regP\[26\] _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4846_ _1036_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _0891_ _0910_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3744__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ _2676_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4941__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3728_ dacArea_dac_cnt_4\[3\] net29 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6447_ _2620_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3483__I _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3659_ _3177_ _3188_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6694__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6378_ _2542_ _2553_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5329_ _1509_ _1510_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5249__A2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A3 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6685__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3499__A1 dspArea_regP\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3499__B2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5822__B _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4160__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4999__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _0834_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _1862_ _1863_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _0815_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4923__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _0746_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _2458_ _2474_ _2477_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3513_ _3077_ _3078_ net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4493_ _0628_ _0685_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6232_ _2324_ _2325_ _2322_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3444_ dspArea_regP\[36\] _2992_ _3006_ _3021_ _3022_ dspArea_regP\[4\] _3023_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6163_ _2161_ _2260_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _1288_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _2133_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_57_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5100__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _1134_ _1136_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_66_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5651__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3414__A1 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5947_ _0195_ dspArea_regA\[20\] _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3478__I _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5878_ _2022_ _2054_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I wb_ADR[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5167__A1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4829_ _1019_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4390__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6825__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5945__A3 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4133__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3892__A1 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3644__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _0004_ net65 dacArea_dac_cnt_4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1981_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5397__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ dspArea_regP\[40\] _2942_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _0207_ net122 _0170_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5732_ _1894_ _1896_ _1913_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5663_ _1844_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4614_ _0755_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _1669_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4545_ _0736_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6649__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4476_ _0596_ _0598_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6215_ _2297_ _2298_ _2295_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4124__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ _3008_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6848__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _2219_ _2249_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _2096_ _2255_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _1210_ _1211_ _1216_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3635__A1 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input10_I la_data_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5312__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6812__A1 dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5615__A2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3626__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6040__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4354__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4330_ _0172_ _3037_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5303__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _0406_ _3015_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6000_ _0242_ _3050_ _2092_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5854__A2 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _0347_ _0350_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input2_I la_data_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6902_ _0056_ clknet_3_5__leaf_wb_clk_i dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6833_ _0141_ net65 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _2843_ _2880_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4042__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3976_ _0193_ net119 _0170_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5715_ _1823_ _1897_ _1832_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6695_ _2824_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5646_ _1826_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5542__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5577_ _1571_ _1760_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_2_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4528_ _0223_ _3001_ _0643_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I la_data_in[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4459_ _0404_ _3020_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3856__A1 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _0232_ _3066_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5781__A1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4887__A3 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5836__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3847__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6261__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4272__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3830_ _3321_ _3320_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_32_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3761_ _3265_ _3267_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4575__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ _1605_ _1608_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6480_ _2584_ _2585_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3692_ dacArea_dac_cnt_3\[3\] net20 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _0183_ _3081_ _1425_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _1547_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _0203_ _3009_ _0461_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XDSP48_208 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_219 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5293_ _1471_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7032_ net144 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5827__A2 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _0437_ _0439_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4175_ dspArea_regP\[5\] _0168_ _3025_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_28_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input112_I wb_DAT_MOSI[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _3111_ _2975_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_24_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _0244_ _3106_ _2859_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_52_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3959_ _0166_ _0179_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_17_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6678_ dspArea_regP\[37\] _0259_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5629_ _0212_ _3061_ _1603_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4318__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5515__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6243__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4780__I _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4309__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6909__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _2157_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4931_ _1114_ _1115_ _1120_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4796__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _0792_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _2730_ _2731_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3813_ _3308_ _3306_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4793_ _0914_ _0984_ _0923_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6532_ dspArea_regP\[33\] _2667_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3744_ dacArea_dac_cnt_4\[6\] net32 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6463_ _2337_ _2340_ _2633_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3675_ dacArea_dac_cnt_3\[0\] net17 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5414_ _1596_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _2499_ _0297_ _2569_ _1461_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xoutput133 net133 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput144 net144 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _1524_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput155 net155 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput166 net166 wb_DAT_MISO[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput177 net177 wb_DAT_MISO[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput188 net188 wb_DAT_MISO[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5276_ _1371_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7015_ net143 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6473__A2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ _0375_ _0425_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4484__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4158_ _0190_ _3008_ _0334_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _0273_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3444__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5984__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__I _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3944__I dspArea_regB\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4475__A1 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4015__I _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput13 la_data_in[20] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 la_data_in[30] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput35 la_data_in[40] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 la_data_in[50] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput57 la_data_in[60] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput68 wb_ADR[11] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput79 wb_ADR[21] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5274__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ _3035_ net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _1317_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6455__A2 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5061_ _1167_ _1247_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__6881__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4466__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _0223_ net101 _0169_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4218__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ _2142_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5966__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _1103_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ _1978_ _0297_ _2075_ _1461_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_61_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5718__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4845_ _0925_ _0942_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_32_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _0895_ _0909_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_14_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _2681_ _2688_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3727_ _3234_ _3241_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4941__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _2542_ _2553_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3658_ dacArea_dac_cnt_2\[4\] net13 _3187_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__6694__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ _2545_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3589_ _3118_ _3133_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _1511_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input40_I la_data_in[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _1443_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6134__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6685__A2 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3499__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4620__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _0820_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6373__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4561_ _0750_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4923__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _2475_ _2407_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3512_ dspArea_regP\[17\] _3072_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3982__I0 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6125__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _0578_ _0686_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6231_ _2324_ _2325_ _2322_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6676__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3443_ _3003_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _1964_ _2070_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5113_ _1293_ _1298_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _2123_ _2134_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _1134_ _1136_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5100__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _0404_ _3085_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5877_ _2057_ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _0176_ _3056_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input88_I wb_ADR[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _0863_ _0866_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_4_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _2602_ _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3892__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _1879_ _1891_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6780_ _3111_ _2946_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _0206_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5397__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5731_ _1894_ _1896_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ _1727_ _1729_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _0805_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5593_ _1672_ _1680_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4544_ _0737_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_7_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ dspArea_regP\[10\] _0597_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _2297_ _2298_ _2295_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3426_ _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _2323_ _2248_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _2149_ _2152_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5085__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _1210_ _1211_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3635__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4832__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3399__A1 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _0205_ _3079_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_16_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__I _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5312__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3874__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6942__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4023__I _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _0201_ _3008_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5303__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4191_ _0357_ _0388_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3865__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__B _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__B2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3617__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6901_ _0055_ clknet_3_6__leaf_wb_clk_i dspArea_regA\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _0140_ net65 dacArea_dac_cnt_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _2904_ _2926_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3975_ _0192_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4042__A2 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ _1824_ _1825_ _1830_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6694_ _0244_ _3094_ _2825_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _1827_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5576_ _1574_ _1756_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5542__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _0639_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4458_ _0593_ _0651_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6965__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3409_ _2991_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4389_ _0201_ _3016_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3856__A2 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _2305_ _2306_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _2236_ _2237_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5648__B _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3947__I _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6323__I dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A2 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6730__A1 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5533__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3544__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5836__A3 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5049__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6797__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4272__A2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4018__I _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5221__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3760_ dacArea_dac_cnt_5\[2\] net37 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__A1 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3691_ dacArea_dac_cnt_3\[3\] net20 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_12_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5430_ _1614_ _1615_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6721__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _1384_ _1447_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4312_ _0407_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5292_ _1477_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XDSP48_209 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5288__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7031_ net143 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4243_ _0355_ _0442_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3838__A2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5460__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input105_I wb_DAT_MOSI[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ dspArea_regP\[47\] _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6746_ _2889_ _2893_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3958_ _0178_ net116 _0170_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3774__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6677_ _0299_ _2846_ _2847_ _1461_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3889_ _3038_ _3360_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6712__A1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _1808_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5515__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input70_I wb_ADR[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _1706_ _1739_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A1 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A2 dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5506__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3517__A1 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5442__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4930_ _1114_ _1115_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4861_ _1048_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6600_ _2771_ _2729_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ dacArea_dac_cnt_6\[5\] net49 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5745__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _0915_ _0916_ _0921_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3743_ _3234_ _3254_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6531_ _2645_ _0297_ _2704_ _1461_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3674_ _3112_ _3200_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6462_ _2564_ _2635_ _2636_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _1597_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6393_ _0792_ _2567_ _2568_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_12_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput134 net134 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_47_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ _1528_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xoutput145 net145 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput156 net156 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput167 net167 wb_DAT_MISO[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput178 net178 wb_DAT_MISO[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput189 net189 wb_DAT_MISO[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5275_ _1374_ _1382_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _0378_ _0382_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4157_ _0184_ _3017_ _0300_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4088_ _0287_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_3_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5433__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__C2 dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3497__I _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3747__A1 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _2896_ _2897_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6464__A3 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 la_data_in[21] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput25 la_data_in[31] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 la_data_in[41] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput47 la_data_in[51] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput58 la_data_in[61] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput69 wb_ADR[12] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _1086_ _1248_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ _0222_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4466__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _2041_ _2047_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _0634_ _3025_ _0994_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5893_ _1773_ _2074_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4206__I _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5718__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4844_ _0938_ _0941_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _0884_ _0885_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6514_ _2686_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3726_ dacArea_dac_cnt_4\[3\] net29 _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6445_ _2545_ _2552_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3657_ _3185_ _3183_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6376_ _2550_ _2551_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3588_ dacArea_dac_cnt_0\[5\] net56 _3132_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5327_ _1512_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_57_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _1306_ _1444_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input33_I la_data_in[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ _0405_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5189_ _0236_ _3026_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5406__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5957__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__I dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6134__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5893__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6918__D _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4448__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5948__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4620__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6373__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4560_ _0751_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_15_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3511_ _3076_ _2999_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3982__I1 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4491_ _0608_ _0609_ _0607_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_7_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4136__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3442_ _3020_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6230_ _2391_ _2394_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _2338_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _1299_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1226_ _1230_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6061__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5945_ _0188_ _3093_ _2040_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_43_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3976__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _1930_ _1946_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _0180_ _3052_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _0887_ _0947_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3709_ net146 net25 _3227_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4689_ _0729_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6428_ _2517_ _2532_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6359_ _2429_ _2431_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6871__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5866__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5618__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _0205_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5730_ _1898_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5661_ dspArea_regP\[22\] _1728_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4612_ _0731_ _0740_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5592_ _1667_ _1774_ _1775_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _0218_ _3007_ _0638_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3580__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6649__A3 _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _0667_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5857__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3425_ dspArea_regA\[1\] _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _2245_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _2149_ _2152_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5085__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5026_ _1212_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_2_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4832__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6034__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4596__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6894__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ _0209_ _3074_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5859_ _2037_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3901__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5895__I dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6328__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4304__I _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4339__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4190_ _0330_ _0389_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_45_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6167__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _0054_ clknet_3_6__leaf_wb_clk_i dspArea_regA\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _0139_ net65 dacArea_dac_cnt_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6762_ _2910_ _0297_ _2929_ _3109_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3974_ dspArea_regB\[5\] _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5713_ _1807_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6693_ _2861_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6319__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A3 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ _0193_ _3080_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5575_ _1574_ _1756_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3553__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4526_ _0642_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4750__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4457_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4502__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3408_ net91 _2986_ _2990_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4388_ _0583_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _2235_ _2243_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _0178_ _3105_ _2124_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4805__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5009_ _0212_ _3037_ _0993_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3963__I _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3544__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__A1 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__A1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5297__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5221__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5772__A3 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4034__I _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3783__A2 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _3177_ _3212_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _1443_ _1446_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4311_ _0196_ _3015_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ _0241_ _3026_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6485__A1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ net151 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4242_ dspArea_regP\[7\] _0440_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _0370_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6788__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _3142_ _2973_ _2974_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_1_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6745_ _2844_ _2905_ _2904_ _2912_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3957_ _0177_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_32_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4971__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ dspArea_regP\[36\] _0874_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3888_ net122 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6932__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5627_ _1809_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4723__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _1741_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input63_I la_data_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _0559_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5489_ _0972_ _3038_ _1599_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6476__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5279__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__C _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6334__I _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5203__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3517__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6467__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4493__A3 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4029__I _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4860_ _1050_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3811_ _3292_ _3307_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6955__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _0899_ _0908_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6530_ _0792_ _2702_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3742_ dacArea_dac_cnt_4\[6\] net32 _3253_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6461_ _2501_ _2563_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3673_ net145 net16 _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4705__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ _0222_ _3044_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6392_ _2501_ _2503_ _2566_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _1429_ _1431_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xoutput135 net135 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput146 net146 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput157 net157 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput168 net168 wb_DAT_MISO[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput179 net179 wb_DAT_MISO[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _0792_ _1459_ _1460_ _1461_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4225_ _0378_ _0382_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5681__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4156_ _0325_ _0326_ _0328_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_28_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ _0289_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6630__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5433__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3444__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__B2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4989_ _0241_ _3013_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _2858_ _2866_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__3747__A2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__A1 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6659_ _2815_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5121__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5424__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5727__A3 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3738__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4935__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput15 la_data_in[22] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput26 la_data_in[32] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 la_data_in[42] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput48 la_data_in[52] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput59 la_data_in[62] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3910__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ _0221_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3674__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5415__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _2043_ _2046_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _0212_ _3033_ _0902_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5892_ _2070_ _2073_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _1017_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_18_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4423__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4926__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4774_ _0880_ _0886_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_18_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _0242_ _3081_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3725_ dacArea_dac_cnt_4\[2\] net28 _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6444_ _2614_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3656_ dacArea_dac_cnt_2\[3\] net11 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5351__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _0241_ _3070_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3587_ _3130_ _3131_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ _0406_ _3065_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3901__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _1339_ _1340_ _1338_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4208_ _0365_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_5_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _0233_ _3026_ _1292_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA_input26_I la_data_in[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4139_ dspArea_regP\[4\] _0306_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5406__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5342__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__I _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5893__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3904__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3408__A1 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4908__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3510_ _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _0608_ _0609_ _0607_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4136__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3441_ _3019_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5333__A1 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__A2 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _2176_ _2259_ _2157_ _2160_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5111_ _0634_ _3034_ _1197_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _2191_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5042_ _1131_ _1133_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6061__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5944_ _1933_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4072__A1 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ _1942_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _0186_ _3048_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _0827_ _0948_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ _3225_ _3223_ _3226_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6116__A3 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4688_ _0226_ _3011_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _2518_ _2531_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4127__A2 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3639_ _3142_ _3171_ _3172_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6358_ _2513_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3886__A1 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _1494_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6289_ _0228_ _3081_ _2310_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6052__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__A1 dspArea_regP\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6043__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ dspArea_regB\[8\] _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3801__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _1841_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4611_ _0736_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5591_ _1752_ _1753_ _1749_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4542_ _0212_ _3016_ _0573_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5306__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ dspArea_regP\[11\] _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6212_ _2367_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5857__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3424_ _2998_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _2295_ _2299_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5609__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _2196_ _2250_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _1213_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4293__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A1 dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5927_ _0216_ _3069_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _2038_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I wb_ADR[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5545__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _0982_ _0983_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_6_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _1159_ _1252_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5848__A2 dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4520__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6273__A2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__A2 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4339__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__I0 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6830_ _0138_ net65 dacArea_dac_cnt_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _0874_ _2927_ _2928_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3973_ _0166_ _0191_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _1812_ _1815_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_17_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _0243_ _3098_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5790__A4 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ _0196_ _3075_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5527__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5574_ _1755_ _1758_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4525_ _0717_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _0182_ _0178_ _3037_ _3033_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3407_ net88 _2989_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _0190_ _3026_ _0525_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_8_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6126_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_59_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6255__A2 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6057_ _2124_ _2139_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6861__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _1194_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3474__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _0113_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6191__A1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4257__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4310_ _0505_ _0506_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_5290_ _1475_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ _0250_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6485__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6884__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4172_ _0371_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4799__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6813_ dspArea_regP\[46\] _0250_ _2966_ _2971_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__5748__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _2878_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3956_ _0176_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _2844_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3887_ _3364_ _3347_ _3365_ _3350_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5626_ _0205_ _3064_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5920__A1 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _1627_ _1644_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4508_ _0698_ _0699_ _0701_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_144_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _0229_ _3046_ _1490_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input56_I la_data_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _0634_ _3008_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_78_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6228__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6109_ _2129_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_59_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5739__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5675__B _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6164__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3907__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A3 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3438__C1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4650__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3810_ dacArea_dac_cnt_6\[5\] net49 _3306_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4790_ _0904_ _0907_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6460_ _2489_ _2491_ _2565_ _2486_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3672_ _3197_ _3195_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5411_ _0226_ _3040_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6391_ _2501_ _2503_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5342_ dspArea_regP\[19\] _1430_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput136 net136 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput147 net147 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput158 net158 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput169 net169 wb_DAT_MISO[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5273_ _3109_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _0417_ _0421_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4155_ _0323_ _0352_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3692__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _0178_ _3002_ _0268_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_55_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input110_I wb_DAT_MOSI[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4641__A1 _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4988_ _1176_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6727_ _2855_ _2857_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_20_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3939_ _0162_ _3348_ _0163_ _0157_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4944__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _2817_ _2828_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _0240_ _3038_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6589_ dspArea_regP\[34\] _2717_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5121__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3969__I _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 la_data_in[23] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 la_data_in[33] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 la_data_in[43] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput49 la_data_in[53] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5360__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3879__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6922__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _2137_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4623__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _1098_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5891_ _2071_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4842_ _1030_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_20_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4926__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ _0877_ _0963_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6512_ _2684_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3724_ _3236_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ dacArea_dac_cnt_2\[3\] net11 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6443_ _2616_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6374_ _2548_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3586_ dacArea_dac_cnt_0\[4\] net45 _3128_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5351__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ _0196_ _3061_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5256_ _1339_ _1340_ _1338_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _0406_ _3011_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _0228_ _3034_ _1191_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_68_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3665__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4862__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _0337_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_29_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input19_I la_data_in[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _0261_ _0270_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3976__I0 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5342__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6945__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3440_ dspArea_regA\[4\] _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6530__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _0213_ _3041_ _1100_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _0243_ _3054_ _2192_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5097__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ dspArea_regP\[16\] _1132_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4993__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _0181_ _3101_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _1944_ _2055_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _1006_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6818__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3958__I0 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5572__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _0860_ _0861_ _0859_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3707_ dacArea_dac_cnt_3\[6\] net24 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _0878_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6426_ _2599_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3638_ dacArea_dac_cnt_2\[0\] net8 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_49_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5324__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6968__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6357_ _2517_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_1_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3569_ _3111_ _3116_ _3117_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3886__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ _0206_ _3052_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _2462_ _2463_ _2464_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _1423_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5012__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5563__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3574__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6512__A1 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3877__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4826__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6579__A1 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4053__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ _0739_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5590_ _1752_ _1753_ _1749_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_15_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3565__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4541_ _0732_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5306__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4472_ _0167_ _3049_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3423_ _3005_ net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6211_ _2370_ _2373_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_48_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3868__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _2303_ _2307_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_48_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _2120_ _2251_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_58_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _0406_ _3052_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6282__A3 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5926_ _2103_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__A3 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5857_ _0177_ _3101_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _0985_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5788_ _1967_ _1970_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input86_I wb_ADR[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3556__A1 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _0173_ _3057_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6409_ _2582_ _2583_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3859__A2 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4284__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5784__A2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6584__I1 _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6760_ _2911_ _2913_ _2926_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _0190_ net118 _0170_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5711_ _1812_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6691_ _2859_ _0238_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5642_ _0201_ _3069_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5527__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3538__A1 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ _1574_ _1756_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4524_ _0629_ _0718_ _0717_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4455_ _0582_ _0594_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3406_ _2987_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4386_ _0467_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4502__A3 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3710__A1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _2239_ _2242_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6056_ _2138_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4266__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _1195_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3474__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3474__C2 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _0112_ clknet_3_6__leaf_wb_clk_i dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _2087_ _2088_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6889_ _0043_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3529__A1 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3500__I _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A2 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4331__I dspArea_regB\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _0398_ _0437_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4171_ _0176_ _3019_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ dspArea_regP\[46\] _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3410__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5748__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3759__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6743_ _2900_ _2903_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_23_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3955_ dspArea_regB\[2\] _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _2843_ _2804_ _2809_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3886_ _3034_ _3360_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5625_ _0209_ _3060_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4241__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4184__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5556_ _1639_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5920__A2 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ _0700_ _0553_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5487_ _1671_ _1609_ _1612_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _0217_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5684__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I la_data_in[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4369_ _0211_ _3007_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _0196_ _3097_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _2217_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_46_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6117__B _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6164__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4175__A1 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3922__A1 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__I0 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6219__A3 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__I _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3438__C2 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4650__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _3250_ _3248_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3671_ dacArea_dac_cnt_2\[6\] net15 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _0231_ _3037_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6390_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5341_ _1525_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput137 net137 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput148 net148 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput159 net159 wb_ACK vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5272_ dspArea_regP\[19\] _0874_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4223_ _0379_ _0381_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4154_ _3110_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4085_ _0288_ _0267_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input103_I wb_DAT_MOSI[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4987_ _1173_ _1174_ _1175_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6726_ _2886_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3938_ _3102_ _3383_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6657_ _2819_ _2827_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3869_ net116 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4157__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5608_ _1790_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6588_ _2740_ _2743_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5539_ _1722_ _1723_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5409__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__I _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6874__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 la_data_in[24] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 la_data_in[34] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput39 la_data_in[44] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5896__A1 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5648__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4623__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5820__A1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _1099_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5890_ _1964_ _1975_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_61_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _0931_ _1031_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3895__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4387__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ _0951_ _0953_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _0237_ _3086_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3723_ dacArea_dac_cnt_4\[2\] net28 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4139__A1 dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6442_ _2538_ _2554_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3654_ _3177_ _3184_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6373_ _0237_ _3076_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6220__B _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3585_ dacArea_dac_cnt_0\[4\] net45 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5324_ _0201_ _3057_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5255_ _1408_ _1439_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4311__A1 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _0192_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _1373_ _1302_ _1305_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ dspArea_regP\[5\] _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6064__A1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _0215_ _0272_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_25_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5811__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6897__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__A2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6709_ _2853_ _2854_ _2877_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3976__I1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A1 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6358__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5869__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _1227_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5942_ _2121_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ _1839_ _1847_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _1014_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5021__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3958__I1 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _0860_ _0861_ _0859_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3583__A2 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3706_ dacArea_dac_cnt_3\[6\] net24 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4686_ _0807_ _0826_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6425_ _2550_ _2551_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3637_ dacArea_dac_cnt_2\[0\] net8 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6356_ _2518_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3568_ _3114_ _3115_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_1_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _0210_ _3048_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6287_ _2373_ _2388_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3499_ dspArea_regP\[47\] _2991_ _2998_ _3066_ _3003_ dspArea_regP\[15\] _3067_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5238_ _1424_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_76_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input31_I la_data_in[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__I _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5169_ _1167_ _1351_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_29_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__A2 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5012__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4360__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4299__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_192 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3503__I _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6579__A2 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__B1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _0733_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4762__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4471_ _0174_ _3045_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6210_ _2378_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3422_ dspArea_regP\[32\] _2992_ _2999_ _3002_ _3004_ dspArea_regP\[0\] _3005_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2312_ _2316_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_48_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2146_ _2147_ _2145_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _0196_ _3049_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6019__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5490__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5242__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5925_ _2104_ _2105_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _0181_ _3097_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5784__B _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4807_ _0990_ _0995_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_22_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5787_ _1776_ _1865_ _1966_ _1765_ _1969_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3556__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input79_I wb_ADR[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _0827_ _0859_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5075__I _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _0207_ dspArea_regA\[24\] _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6339_ _2446_ _2448_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4808__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4154__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4992__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4090__S _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3926__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6249__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4329__I _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5224__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6958__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3971_ _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5710_ _1815_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4983__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6690_ _2763_ _2856_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _0190_ _3081_ _1724_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3538__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _1655_ _1658_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _0633_ _0646_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_7_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _0648_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3405_ net93 net95 net94 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _0182_ _3033_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6124_ _2300_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _2233_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5006_ _0205_ _3040_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_61_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5779__B _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3474__A1 dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3474__B2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6412__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6957_ _0111_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3777__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _0236_ _3054_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4974__A1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6888_ _0042_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5839_ _2000_ _2002_ _2019_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3529__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A1 _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6479__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3701__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6651__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3768__A2 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5142__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _0181_ _3015_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6811_ _3142_ _2970_ _2972_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ dspArea_regP\[39\] _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3954_ _0166_ _0175_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4420__A3 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6673_ _2804_ _2809_ _2843_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3885_ net121 _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4708__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5624_ _0216_ _3057_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5555_ _1642_ _1647_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ _0700_ _0553_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _1517_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5133__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4437_ _0631_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4368_ _0506_ _0507_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3695__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6107_ _2232_ _2241_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0299_ _0496_ _0497_ _0157_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__A1 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _2198_ _2200_ _2216_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4947__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4432__I _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4175__A2 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3922__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__I1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5124__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3438__A1 dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3438__B2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ dacArea_dac_cnt_2\[6\] net15 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5363__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ dspArea_regP\[20\] _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput127 net127 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput138 net138 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput149 net149 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_5_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5271_ _1454_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6458__A4 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4222_ dspArea_regP\[6\] _0380_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5666__A2 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3677__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4153_ _0299_ _0353_ _0354_ _0157_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_28_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _0265_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3421__I _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4986_ _1173_ _1174_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6725_ _2889_ _2893_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3937_ net114 _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _2825_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3868_ _3351_ _3347_ _3352_ _3350_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _1787_ _1788_ _1789_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4157__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _2735_ _2739_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3799_ dacArea_dac_cnt_6\[2\] net46 _3297_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3904__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5538_ dspArea_regB\[2\] dspArea_regA\[20\] _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input61_I la_data_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5106__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _1589_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output148_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6606__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 la_data_in[25] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 la_data_in[35] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5345__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3659__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ _0935_ _0937_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4387__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _0951_ _0953_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6510_ _2682_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3722_ _3234_ _3237_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6441_ _2615_ _2537_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3653_ dacArea_dac_cnt_2\[3\] net11 _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_9_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _2546_ _2547_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3584_ _3118_ _3129_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5323_ _0190_ _3066_ _1426_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__3416__I _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5254_ _1440_ _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_9_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ _0404_ _3000_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4311__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ _1218_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _0167_ _3025_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4247__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4067_ dspArea_regP\[2\] _0271_ _0259_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4378__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5575__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _1066_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6708_ _2853_ _2854_ _2877_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ dspArea_regP\[35\] _2768_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3889__A1 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4302__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5541__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6841__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3996__I _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6547__I _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6294__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4057__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _0202_ _3081_ _2031_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_80_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ _2036_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_21_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _1007_ _1008_ _1013_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4754_ _0911_ _0943_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3705_ _3177_ _3224_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4685_ _0811_ _0825_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__4530__I _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3636_ _3112_ _3170_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6424_ _2598_ _2549_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6355_ _2523_ _2528_ _2530_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3567_ _3114_ _3115_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6809__A1 dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _0218_ _3045_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6286_ _2373_ _2388_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3498_ _3065_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5237_ dspArea_regB\[2\] _3074_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6864__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _1155_ _1158_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input24_I la_data_in[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ _0299_ _0320_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ _1209_ _1287_ _1218_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5012__A3 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4220__A1 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6276__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XDSP48_193 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6028__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5787__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__A3 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4514__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5711__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _2317_ _2318_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A2 dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _2146_ _2147_ _2145_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4278__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _0201_ _3045_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6019__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ dspArea_regB\[11\] _3064_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_53_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5855_ _0188_ _3093_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ _0996_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5784__C _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4202__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _1867_ _1968_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4737_ _0926_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4668_ _0860_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3619_ _3155_ _3153_ _3156_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6407_ _0211_ _3101_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5702__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _0711_ _0786_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _2441_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6269_ _2442_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6430__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5941__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3942__C _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6249__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ _0188_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _0184_ _3090_ _1630_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_31_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5571_ _1655_ _1658_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5932__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4522_ _0633_ _0646_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4453_ _0203_ _3016_ _0589_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3404_ net92 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4384_ _0579_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _2206_ _2301_ _2300_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3424__I _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _0202_ _3086_ _2130_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__3459__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5005_ _0209_ _3036_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_38_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3474__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input126_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6902__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _0110_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _0233_ _3054_ _2008_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _0041_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6176__A1 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ _2000_ _2002_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_14_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input91_I wb_ADR[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5923__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _1854_ _1855_ _1853_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_33_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output178_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6651__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6380__I _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4717__A2 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3509__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5142__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6925__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6810_ _0298_ _2958_ _2963_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _0299_ _2908_ _2909_ _3109_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3953_ _0174_ net110 _0170_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6158__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6672_ _2838_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3884_ _3362_ _3347_ _3363_ _3350_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _1803_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3419__I _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5554_ _1720_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4505_ _0549_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5485_ _1508_ _1518_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4436_ _0581_ _0591_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5133__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _0562_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ dspArea_regP\[28\] _2223_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ dspArea_regP\[8\] _0299_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6633__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _2198_ _2200_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ _0093_ clknet_3_7__leaf_wb_clk_i dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4947__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4175__A3 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3999__I _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3438__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput128 net128 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput139 net139 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_5270_ _1455_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ _0418_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4874__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4152_ dspArea_regP\[5\] _0299_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__I _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6615__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4083_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4985_ _0237_ _3017_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3988__I0 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6724_ _2890_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3936_ _0160_ _3348_ _0161_ _0157_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3601__A2 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6655_ _0243_ _3094_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _3009_ _3348_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5606_ _1787_ _1788_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5354__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ dspArea_regP\[35\] _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3798_ _3294_ _3296_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5537_ _0180_ _3084_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _1651_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input54_I la_data_in[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4419_ _0568_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3668__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5399_ _1583_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6606__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4871__C _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5593__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 la_data_in[26] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3522__I _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6781__A1 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ dspArea_regP\[15\] _0259_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5584__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ dacArea_dac_cnt_4\[2\] net28 _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_18_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _2534_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3652_ dacArea_dac_cnt_2\[2\] net10 _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6533__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3583_ dacArea_dac_cnt_0\[4\] net45 _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_6371_ _0972_ _3076_ _2440_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3898__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ _0184_ _3076_ _1323_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _1320_ _1337_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _0200_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5184_ _1209_ _1219_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_68_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _0174_ _3020_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3432__I _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _0261_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_83_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5272__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5024__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _1155_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ _2872_ _2876_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3919_ _3076_ _3383_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4899_ _0990_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _2805_ _2806_ _2808_ _2796_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_22_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6569_ _2676_ _2689_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5094__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3889__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4438__I _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4057__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _0198_ _3090_ _1924_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5871_ _2048_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5006__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _1007_ _1008_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4753_ _0944_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ dacArea_dac_cnt_3\[6\] net24 _3223_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6506__A1 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ _0644_ _0798_ _0802_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_6423_ _2548_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3635_ net144 net7 _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__3427__I _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6354_ _2442_ _2445_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3566_ dacArea_dac_cnt_0\[1\] net12 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6809__A2 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _1488_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6285_ _2370_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3497_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5236_ _0180_ _3068_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5167_ _1070_ _1154_ _1251_ _1163_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4118_ _0316_ _0319_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _1210_ _1211_ _1216_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4048__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__A1 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I la_data_in[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4049_ dspArea_regP\[1\] _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5817__I _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__S _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_194 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_47_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__A1 _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5787__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _2993_ net91 _2986_ _2989_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_48_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3722__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _2219_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4278__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I la_data_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5021_ _0190_ _3054_ _1128_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5227__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5923_ _0225_ _3060_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5854_ _2025_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_80_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4805_ _0218_ _3020_ _0903_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_10_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5785_ _1776_ _1865_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4202__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4736_ _0927_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5950__A2 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4667_ _0757_ _0773_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6831__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ _2577_ _2580_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3618_ dacArea_dac_cnt_1\[3\] net3 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5702__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3713__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6337_ _2508_ _2512_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3549_ dspArea_regP\[24\] _3004_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6268_ _2443_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4269__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5219_ _1386_ _1388_ _1405_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6199_ _2375_ _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_40_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5218__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4441__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6718__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__B _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5209__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6185__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6854__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _1667_ _1749_ _1754_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__5932__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _0628_ _0714_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_144_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4452_ _0198_ _3026_ _0517_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4499__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3403_ _2982_ _2985_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4383_ _0203_ _3013_ _0518_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _2212_ _2213_ _2211_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _2030_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_39_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3459__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3459__C2 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5004_ _0216_ _3033_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input119_I wb_DAT_MOSI[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _0109_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5906_ _0228_ _3062_ _1901_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _0040_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ _2004_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6176__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ _1916_ _1947_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input84_I wb_ADR[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4719_ _0197_ _3038_ _0753_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5699_ _1881_ _1816_ _1819_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5439__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5611__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6877__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5914__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3925__A1 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ dspArea_regP\[38\] _0299_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _0173_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_56_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6671_ _2839_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3883_ _3030_ _3360_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4169__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _1804_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3916__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5553_ _1733_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4504_ _0499_ _0491_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5484_ _1584_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5669__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _0630_ _0590_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4341__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4366_ _0501_ _0548_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6469__I0 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _2271_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _0445_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2202_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5841__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _0092_ clknet_3_2__leaf_wb_clk_i dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _0023_ net65 dacArea_dac_cnt_6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output190_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4580__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4399__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput129 net129 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ dspArea_regP\[7\] _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _0323_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_68_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _0280_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5823__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _0972_ _3017_ _1096_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6723_ _2891_ _2862_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3935_ _3098_ _3383_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3988__I1 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6654_ _2823_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3866_ net110 _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6000__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ _0236_ _3042_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6585_ _3111_ _2757_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3797_ dacArea_dac_cnt_6\[2\] net46 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5536_ _0186_ _3080_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5467_ _1505_ _1541_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4418_ _0611_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5398_ _1580_ _1581_ _1582_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input47_I la_data_in[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4349_ _0451_ _0486_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6019_ _2112_ _2115_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6058__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6781__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _3235_ _3233_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3595__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _3179_ _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6533__A2 _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _0228_ _3086_ _2376_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3582_ _3126_ _3124_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _1506_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5252_ _1333_ _1336_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ _0401_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5183_ _1277_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ _0268_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_37_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input101_I wb_DAT_MOSI[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6221__A1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4967_ _0880_ _0886_ _1156_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_33_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6706_ _2873_ _2875_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3918_ net107 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3586__A2 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4898_ _0995_ _0998_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_32_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6637_ _2799_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3849_ _3336_ _3334_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4535__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ _2681_ _2688_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5519_ _1684_ _1686_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _2607_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4838__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3577__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4774__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6451__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _2049_ _2050_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6203__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4821_ _1009_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _0841_ _0858_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ dacArea_dac_cnt_3\[5\] net22 _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4683_ _0868_ _0870_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6422_ _2593_ _2596_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3634_ _3167_ _3165_ _3168_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _0207_ _3098_ _2443_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3565_ _3112_ _3113_ _3114_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5304_ _1489_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3871__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6284_ _2459_ _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3496_ dspArea_regA\[15\] _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5235_ _0186_ _3065_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3443__I _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6690__A1 _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _1159_ _1252_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ _0316_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5097_ _1193_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _0168_ _3009_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_71_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _2177_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5548__A3 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3731__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5054__B _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6681__A1 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_195 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6433__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5236__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4278__A3 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _0184_ _3062_ _1020_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5227__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A3 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__I _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ dspArea_regB\[13\] _3057_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5853_ _2033_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4804_ _0211_ _3029_ _0818_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_21_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5784_ _1558_ _1559_ _1767_ _1966_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_21_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4735_ _0176_ _3052_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4666_ _0769_ _0772_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _2578_ _2579_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3617_ dacArea_dac_cnt_1\[3\] net3 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4597_ _0248_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6336_ dspArea_regP\[31\] _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_143_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3548_ _3106_ _2999_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _0207_ dspArea_regA\[22\] _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3479_ dspArea_regP\[43\] _2991_ _2998_ _3050_ _3022_ dspArea_regP\[11\] _3051_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5466__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _1386_ _1388_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_9_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _0223_ _3080_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5149_ _1320_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5218__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6718__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__A3 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5991__C _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3704__A2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _0685_ _0688_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _0629_ _0633_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ net77 net66 _2983_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4382_ _0198_ _3021_ _0460_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _2212_ _2213_ _2211_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _0195_ dspArea_regA\[21\] _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3459__A1 dspArea_regP\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3459__B2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _1189_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_79_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4120__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _0108_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5620__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5905_ _2085_ _2018_ _2021_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3631__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _0039_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5836_ _2009_ _2014_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _1948_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4718_ _0891_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5698_ _1718_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input77_I wb_ADR[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4649_ _0181_ _3044_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _2492_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5439__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3870__A1 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5611__A2 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4178__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3925__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5850__A2 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6821__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3951_ _0172_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4372__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6670_ _2840_ _2793_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3882_ net120 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ _0221_ _3052_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__A2 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5366__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3916__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5552_ _1734_ _1735_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4503_ _0445_ _0495_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5118__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _0244_ _3030_ _1585_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4434_ _0585_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4365_ _0545_ _0547_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _2274_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _0491_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2206_ _2211_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5841__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3852__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6937_ _0091_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6868_ _0022_ net65 dacArea_dac_cnt_6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _1908_ _1911_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6799_ _3111_ _2962_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3907__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6002__I _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A2 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__I dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5520__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _0324_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4081_ _0281_ _0282_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _0229_ _3026_ _0988_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_23_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _2861_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3934_ net113 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5339__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _2820_ _2821_ _2822_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3865_ _3344_ _3347_ _3349_ _3350_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_31_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3874__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _0233_ _3042_ _1692_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3796_ _3292_ _3295_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6584_ dspArea_regP\[34\] _2756_ _0874_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _1709_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_30_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _1537_ _1540_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4417_ _0508_ _0612_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5511__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _1580_ _1581_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__6867__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4348_ _0482_ _0485_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4279_ _0421_ _0423_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6018_ _2112_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_74_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6160__C _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__A2 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5750__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3650_ dacArea_dac_cnt_2\[2\] net10 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ dacArea_dac_cnt_0\[3\] net34 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5741__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5320_ _0203_ _3054_ _1417_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_6_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _1422_ _1435_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4202_ _0189_ _3012_ _0373_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _0243_ _3017_ _1278_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_3_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _0331_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _0178_ _3002_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _1043_ _1046_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6705_ _2874_ _2828_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3917_ _3385_ _3371_ _3386_ _3373_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_32_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__I _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0995_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _2795_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3848_ dacArea_dac_cnt_7\[5\] net58 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4535__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _2735_ _2739_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3779_ _3234_ _3282_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_3_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _1688_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6498_ _2668_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5449_ dspArea_regP\[21\] _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4299__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4838__A3 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output146_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5799__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4471__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6212__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5971__A1 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7021__I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6203__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _1010_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3422__C1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5962__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _0854_ _0857_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_18_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3702_ _3221_ _3219_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4682_ _0792_ _0873_ _0875_ _0157_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3633_ dacArea_dac_cnt_1\[6\] net6 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6421_ _2594_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5714__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3564_ dacArea_dac_cnt_0\[0\] net1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6352_ _2524_ _2527_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5303_ _0222_ _3040_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6283_ _0244_ _3062_ _2403_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3495_ _3063_ net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _1411_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3489__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5165_ _1350_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_5_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4116_ _0317_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _1198_ _1201_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6905__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4047_ dspArea_regP\[0\] _0168_ _3002_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4453__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5998_ _2083_ _2095_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4949_ _1023_ _1138_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ _2725_ _2732_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5705__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6130__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4692__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_196 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6433__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4444__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6197__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5944__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7016__I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6121__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6928__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4683__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _0124_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _2025_ _2101_ _2034_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5852_ _2026_ _2027_ _2032_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _0991_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5935__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _1759_ _1866_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4734_ _0180_ _3048_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _0841_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _0222_ _3093_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3616_ _3118_ _3154_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4596_ net125 _2987_ _0246_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_31_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5155__B _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6335_ _2509_ _2510_ _2355_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3547_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6112__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ _0211_ dspArea_regA\[21\] _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3478_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5217_ _1390_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6197_ _0227_ _3075_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _1333_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_input22_I la_data_in[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5079_ _1177_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3401__A2 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5090__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4450_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5145__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3401_ net97 net96 net68 net67 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4381_ _0572_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6120_ _2297_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2227_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3459__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _1190_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_38_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6953_ _0107_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _1928_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3877__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6884_ _0038_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5908__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5835_ _2015_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6581__A1 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _1834_ _1852_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5384__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4717_ _0895_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5697_ _1709_ _1719_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ _0188_ _3041_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _0757_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6318_ _2337_ _2340_ _2343_ _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6249_ _0193_ _3105_ _2355_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__3912__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3870__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3689__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ dspArea_regB\[1\] _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_56_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4810__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3881_ _3359_ _3347_ _3361_ _3350_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_31_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _0225_ _3048_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5366__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _1636_ _1638_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _3173_ _0621_ _0697_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5118__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5482_ _1664_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _0567_ _0576_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4364_ _0551_ _0549_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _2280_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _0399_ _0492_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _2212_ _2213_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input124_I wb_STB vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _0090_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6867_ _0021_ net65 dacArea_dac_cnt_6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ _1908_ _1999_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6798_ dspArea_regP\[43\] _2961_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_13_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5749_ _0180_ dspArea_regA\[21\] _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output176_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5045__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5520__A2 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7024__I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _0269_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _1171_ _1106_ _1109_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_45_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3598__A1 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6721_ _0238_ _2860_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3933_ _0158_ _3348_ _0159_ _0157_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6652_ _2820_ _2821_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5339__A2 dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ _3109_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6531__C _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _0228_ _3050_ _1598_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6583_ _2748_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3795_ dacArea_dac_cnt_6\[2\] net46 _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_30_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5534_ _1717_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _1613_ _1645_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3890__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4416_ _0542_ _0543_ _0541_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5511__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5396_ _0237_ _3034_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4347_ _0508_ _0541_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__3462__I _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4278_ _0470_ _0474_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4078__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6773__I _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2115_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5027__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A2 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _0073_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6527__A1 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A2 dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__A3 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5502__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6058__A3 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5266__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3547__I _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7019__I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ dacArea_dac_cnt_0\[3\] net34 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5741__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _1326_ _1436_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3504__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4201_ _0183_ _3021_ _0333_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5181_ _1367_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _0332_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4063_ _0265_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3807__A2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5009__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4965_ _1043_ _1046_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6704_ _2817_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6509__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _3070_ _3383_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5980__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ _0998_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _2748_ _2797_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3847_ _3292_ _3335_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3457__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _2737_ _2738_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3778_ dacArea_dac_cnt_5\[6\] net41 _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__3743__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _1693_ _1698_ _1701_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_6497_ _2669_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5448_ _0529_ dspArea_regA\[21\] _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input52_I la_data_in[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4299__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5379_ dspArea_regP\[20\] _1565_ _0441_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5248__A1 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4471__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6748__A1 dspArea_regP\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4214__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5411__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6857__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0925_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_18_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3422__B1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3422__C2 dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3701_ dacArea_dac_cnt_3\[5\] net22 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3973__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ dspArea_regP\[13\] _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_18_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _2513_ _2533_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3632_ dacArea_dac_cnt_1\[6\] net6 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5714__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6351_ _2525_ _2526_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3563_ dacArea_dac_cnt_0\[0\] net1 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5302_ _0226_ _3036_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6282_ _0238_ _3066_ _2401_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3494_ dspArea_regP\[46\] _2991_ _2998_ _3062_ _3003_ dspArea_regP\[14\] _3063_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _1419_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3489__B1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3489__C2 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5164_ _1167_ _1351_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4115_ _0273_ _0292_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _1198_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _0215_ _0252_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5650__A1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4453__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _2086_ _2094_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4205__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _1027_ _1029_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _1067_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _2788_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6549_ _2686_ _2687_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4012__S _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6130__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_197 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_21_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4444__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5641__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6197__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4380__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3560__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7032__I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5920_ _2026_ _2027_ _2032_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _2026_ _2027_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__6188__A2 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _0992_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5782_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5935__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4733_ _0187_ _3045_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4664_ _0854_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6403_ _0227_ _3089_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3615_ dacArea_dac_cnt_1\[3\] net3 _3153_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4595_ _2982_ _2988_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6334_ _3106_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3546_ dspArea_regA\[24\] _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6265_ _0218_ _3089_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3477_ _3048_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4123__A1 _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _1395_ _1400_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_6196_ _0232_ _3070_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3470__I _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5147_ _1226_ _1334_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _0242_ _3013_ _1178_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I la_data_in[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A1 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4007__S _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__A3 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A1 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5614__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3928__A1 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7027__I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ net70 net69 net72 net71 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_4380_ _0567_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_4_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _2228_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I la_data_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5001_ _0221_ _3028_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _0106_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _1919_ _1929_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_81_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6883_ _0037_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _0634_ _3061_ _1907_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5908__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3919__A1 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _1848_ _1851_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3893__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _0899_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5696_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4647_ _0830_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3465__I _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4578_ _0769_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3529_ dspArea_regP\[20\] _3004_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__A1 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _2423_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5844__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ _2355_ _2356_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6021__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__B _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6572__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__A1 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A2 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__A1 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3880_ _3026_ _3360_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5550_ _1636_ _1638_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _0297_ _0695_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5481_ _1665_ _1588_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5118__A3 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4326__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4432_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4877__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4363_ _0555_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _0240_ _3058_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _0433_ _0436_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _0634_ _3069_ _2111_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input117_I wb_DAT_MOSI[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0089_ clknet_3_2__leaf_wb_clk_i dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _0020_ net65 dacArea_dac_cnt_6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6003__A1 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ _1911_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6797_ _3142_ _2960_ _2961_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6554__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4565__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _0187_ _3089_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_41_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input82_I wb_ADR[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _1682_ _1748_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output169_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6242__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4308__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5808__A1 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4981_ _1015_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_45_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3598__A2 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _2887_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3932_ _3094_ _3383_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4795__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _0238_ _3098_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3863_ _3002_ _3348_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5602_ _1785_ _1702_ _1705_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _2749_ _2751_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3794_ _3293_ _3291_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5533_ _1710_ _1711_ _1716_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3770__A2 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5464_ _1648_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4415_ _0542_ _0543_ _0541_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5395_ _0972_ _3034_ _1491_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4346_ _0542_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _0418_ _0420_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6016_ _2182_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5275__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6918_ _0072_ clknet_3_7__leaf_wb_clk_i dspArea_regB\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _0003_ net65 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__I0 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4553__A4 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5502__A3 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5266__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5018__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7035__I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4200_ _0360_ _0367_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3504__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _1269_ _1281_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4131_ _0177_ _3016_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _0255_ _0256_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_3_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4768__A1 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _1070_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6703_ _2819_ _2827_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5439__B _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3915_ net106 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ _1073_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3846_ dacArea_dac_cnt_7\[5\] net58 _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6634_ _2630_ _2749_ _2750_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5193__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3777_ dacArea_dac_cnt_5\[5\] net40 _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6565_ _2672_ _2690_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5516_ _1699_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4940__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6496_ _2571_ _2592_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5447_ _0172_ _3089_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3473__I _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5378_ _1555_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input45_I la_data_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4329_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__A2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3734__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5487__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5239__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4998__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3422__A1 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3422__B2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3700_ _3177_ _3220_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4680_ _0250_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_30_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3631_ _3118_ _3166_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5175__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A3 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ _0207_ _3101_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3562_ _3109_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5301_ _0232_ _3033_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ _2452_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3493_ _3061_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5478__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _1412_ _1413_ _1418_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3489__A1 dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3489__B2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5163_ _1247_ _1250_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6427__A1 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ _0287_ _0291_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5094_ _1201_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ dspArea_regP\[0\] _0251_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4989__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2080_ _2174_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_40_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3413__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__I _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4947_ _1027_ _1029_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4878_ _0967_ _1068_ _1067_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_14_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6951__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _2719_ _2734_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5166__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ dacArea_dac_cnt_7\[1\] net53 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _2720_ _2685_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _2587_ _2583_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output151_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4141__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_198 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_47_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5641__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5794__S _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3707__A2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4904__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4380__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__I _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6824__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5850_ _2028_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _0205_ _3032_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5781_ _1960_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5935__A3 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _0914_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5148__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ _0762_ _0855_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3614_ dacArea_dac_cnt_1\[2\] net2 _3152_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6402_ _0232_ _3086_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4594_ _0355_ _0788_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3545_ _3103_ _3104_ net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6333_ _0203_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _2437_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3476_ dspArea_regA\[11\] _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _1401_ _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4123__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _2371_ _2372_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5146_ _1230_ _1232_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5077_ _1263_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_84_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__A3 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4028_ _0236_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _1983_ _2158_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5139__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6639__A1 dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5311__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6847__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A2 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3873__A1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6811__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3928__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A3 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0225_ _3024_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5605__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _0105_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3616__A1 _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5498__I _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6882_ _0036_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5369__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _0212_ _3069_ _1810_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_14_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3919__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _1930_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _0904_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5695_ _1791_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4646_ _0834_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4344__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _0666_ _0770_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6316_ _2334_ _2413_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3528_ _3090_ _2999_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _2421_ _2422_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3459_ dspArea_regP\[39\] _2992_ _3006_ _3034_ _3022_ dspArea_regP\[7\] _3035_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5844__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _0193_ dspArea_regA\[24\] _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_40_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _1310_ _1311_ _1316_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3607__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5357__B _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5532__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__A3 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7038__I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _0626_ _0694_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5480_ _1576_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4431_ _0572_ _0577_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4326__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4362_ _0549_ _0552_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6101_ _2278_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4293_ _0433_ _0436_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _0212_ _3080_ _2012_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3837__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6251__A2 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _0088_ clknet_3_2__leaf_wb_clk_i dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6865_ _0019_ net65 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6003__A2 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1985_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6796_ dspArea_regP\[42\] _0250_ _2958_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5747_ _1919_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4565__A2 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _1744_ _1747_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input75_I wb_ADR[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5514__A1 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0821_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4253__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6902__D _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4308__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4010__I _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _1006_ _1016_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_45_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ net112 _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4795__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _0234_ _3098_ _2765_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3862_ _3346_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_31_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5601_ _1625_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5744__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4547__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _1974_ _2640_ _2753_ _2639_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3793_ dacArea_dac_cnt_6\[1\] net44 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5532_ _1710_ _1711_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5463_ _1519_ _1536_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _0578_ _0607_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_5394_ _0229_ _3042_ _1393_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0464_ _0481_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4276_ dspArea_regP\[7\] _0419_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6908__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2185_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4235__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6917_ _0071_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4786__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6848_ _0002_ net65 dacArea_dac_cnt_3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5735__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ dspArea_regP\[40\] _2945_ _0874_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5586__I1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A1 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5726__A1 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4005__I _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4130_ _0182_ _3012_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__A2 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4061_ dspArea_regP\[1\] _0254_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4768__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _1150_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6702_ _2867_ _2871_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3914_ _3382_ _3371_ _3384_ _3373_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4894_ _1076_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6633_ _1974_ _2640_ _2803_ _2639_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_20_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5717__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3845_ _3332_ _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6564_ _2668_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5193__A2 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3776_ _3279_ _3277_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5515_ _0634_ _3049_ _1604_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ dspArea_regP\[32\] _2570_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4940__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6142__A1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5446_ _1628_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _1558_ _1559_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_4328_ _0522_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input38_I la_data_in[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4259_ _0456_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6880__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A1 dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3929__I _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4447__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3670__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3422__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ dacArea_dac_cnt_1\[6\] net6 _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3561_ net124 net98 _3111_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _1411_ _1486_ _1420_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6280_ _2455_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3492_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5231_ _1412_ _1413_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_143_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3489__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4686__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5162_ _1247_ _1250_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4113_ _0284_ _0311_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _1269_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_68_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4044_ _0168_ _3002_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_49_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4989__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _2154_ _2155_ _2153_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1130_ _1134_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _0970_ _0980_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _2705_ _2718_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3828_ _3173_ _3319_ _3320_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5166__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ _2684_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3759_ _3234_ _3266_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4913__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__I0 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _2650_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _0202_ _3058_ _1514_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4677__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output144_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_199 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A1 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A3 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _0209_ _3028_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A1 _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _1780_ _1961_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6345__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _0766_ _0768_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _2573_ _2574_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3613_ _3149_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ dspArea_regP\[12\] _0787_ _0441_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ dspArea_regP\[30\] _2428_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3544_ dspArea_regP\[23\] _3004_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4371__A3 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6263_ _2438_ _2439_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3475_ _3047_ net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ _0218_ _3037_ _1297_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_69_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6194_ _2289_ _2293_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5320__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5145_ _1230_ _1232_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5076_ _1264_ _1181_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5084__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4027_ dspArea_regB\[14\] _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _2065_ _2068_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _1116_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6336__A1 dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5139__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4898__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5311__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A3 dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A2 dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _0104_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4813__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5901_ _1993_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_47_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6881_ _0035_ net65 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5832_ _2010_ _2013_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5763_ _1942_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4714_ _0905_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6318__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _0242_ _3038_ _1792_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4645_ _0835_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_30_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4576_ _0670_ _0672_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3552__A1 dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _2489_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_143_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6246_ _2421_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3458_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _0196_ _3101_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _1310_ _1311_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA_input20_I la_data_in[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _1146_ _1149_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__C _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3543__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6964__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4638__A4 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3846__A2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__I _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__A1 dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _0624_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__A2 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3534__A1 dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _0355_ _0558_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6100_ _2275_ _2276_ _2277_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4292_ _0487_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__A1 _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _2207_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5039__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _0087_ clknet_3_2__leaf_wb_clk_i dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3958__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6864_ _0018_ net65 dacArea_dac_cnt_5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5815_ _1988_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6795_ dspArea_regP\[42\] _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1927_ _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5677_ _1796_ _1857_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4628_ _0218_ _3012_ _0735_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5514__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input68_I wb_ADR[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3492__I _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4559_ _0752_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5921__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6229_ _2396_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_89_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4253__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5202__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A2 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5505__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A1 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _0155_ _3348_ _0156_ _0157_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ _3346_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_60_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ _1616_ _1626_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6580_ _2752_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3792_ _3110_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5744__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3755__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5531_ _1712_ _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5462_ _1646_ _1647_ _1535_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4413_ _0608_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5393_ _1578_ _1501_ _1504_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4180__A1 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _0477_ _0480_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4275_ _0471_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _2192_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_41_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input122_I wb_DAT_MOSI[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6916_ _0070_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _0001_ net65 dacArea_dac_cnt_3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3487__I _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _2936_ _2944_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5735__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ _1903_ _1908_ _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output174_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__C _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4021__I dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4060_ _0263_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5414__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _0981_ _1151_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_33_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _2868_ _2870_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3913_ _3066_ _3383_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4893_ _1082_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ _2748_ _2752_ _2797_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3844_ dacArea_dac_cnt_7\[4\] net57 _3330_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_32_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5717__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _2671_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3775_ dacArea_dac_cnt_5\[5\] net40 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5514_ _0212_ _3057_ _1495_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6494_ _2645_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5445_ _1629_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4153__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5376_ _1061_ _1065_ _1355_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3900__A1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4327_ _0523_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _0189_ _3016_ _0415_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_41_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__A2 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _0343_ _0346_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3945__I _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5644__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4447__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A2 dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__I _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4383__A1 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ _3110_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3491_ dspArea_regA\[14\] _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4135__A1 _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _1414_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_64_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5161_ _1266_ _1346_ _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_69_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ _0312_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _1272_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _2982_ _2997_ _0247_ _0249_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5994_ _2154_ _2155_ _2153_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6060__A1 _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3949__A1 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4945_ _1024_ _1026_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4876_ _0970_ _0980_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_21_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _2770_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3827_ _3317_ _3318_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6546_ _2705_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3758_ dacArea_dac_cnt_5\[2\] net37 _3265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_14_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6477_ _0634_ _3102_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3972__I1 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3689_ dacArea_dac_cnt_3\[3\] net20 _3211_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4126__A1 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__I0 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _0197_ _3066_ _1416_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA_input50_I la_data_in[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _1481_ _1542_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_47_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5626__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7029_ net150 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__S _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__A1 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5617__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _0915_ _0916_ _0921_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3946__A4 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _0766_ _0768_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6345__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _2528_ _2530_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6870__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3612_ dacArea_dac_cnt_1\[2\] net2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ _0712_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _2478_ _2481_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3543_ _3102_ _2999_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4108__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _0222_ _3085_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3474_ dspArea_regP\[42\] _2991_ _3006_ _3046_ _3022_ dspArea_regP\[10\] _3047_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5856__A1 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _0212_ _3045_ _1196_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6193_ _2224_ _2292_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5144_ _1326_ _1330_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_9_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5075_ _1169_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6281__A1 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _0215_ _0235_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _2065_ _2068_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_12_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3398__A2 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4595__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4928_ _1117_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input98_I wb_CYC vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3495__I _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__A2 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _0955_ _0959_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4898__A2 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _2630_ _2646_ _2701_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5847__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4813__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _0243_ _3046_ _1994_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6880_ _0034_ net65 dacArea_dac_cnt_7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__A1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5831_ _2011_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_62_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ _1840_ _1943_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_61_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4713_ _0217_ _3016_ _0819_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6318__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5693_ _1874_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4204__I _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4644_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4575_ _0670_ _0672_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_11_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3552__A2 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6314_ _2415_ _2416_ _2333_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3526_ dspArea_regA\[20\] _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5829__A1 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _0202_ _3102_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3457_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4501__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _0201_ _3097_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _1312_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ _1146_ _1149_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I la_data_in[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ dspArea_regB\[11\] _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6006__A1 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4568__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5532__A3 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3543__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6245__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6796__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4024__I _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3534__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ dspArea_regP\[9\] _0557_ _0441_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _0360_ _0367_ _0432_ _0489_ _0428_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A1 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _2208_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5287__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I la_data_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5039__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6932_ _0086_ clknet_3_2__leaf_wb_clk_i dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4798__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _0017_ net65 dacArea_dac_cnt_5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _1994_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6794_ _0298_ _2958_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_22_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1920_ _1921_ _1926_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3773__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ _1706_ _1858_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4627_ _0211_ _3020_ _0637_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _0192_ _3032_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3509_ _3074_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4489_ _0647_ _0679_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6228_ _2399_ _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _2176_ _2259_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6931__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6466__A1 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3858__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _2989_ _2996_ _3345_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_32_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ _3173_ _3290_ _3291_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_13_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5530_ _1713_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _1524_ _1531_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4412_ _0521_ _0540_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4704__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _1420_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4343_ _0521_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ dspArea_regP\[8\] _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _0240_ _3054_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6209__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input115_I wb_DAT_MOSI[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6915_ _0069_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _0000_ net65 dacArea_dac_cnt_3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6954__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6777_ _2940_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3989_ _0166_ _0204_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_22_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _1909_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input80_I wb_ADR[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ dspArea_regP\[23\] _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_11_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4934__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6687__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6827__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A1 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4961_ _1039_ _1042_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6700_ _2869_ _2829_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3912_ _3346_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_33_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4892_ _0240_ _3009_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6631_ _2758_ _0297_ _2802_ _1461_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_32_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5178__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3843_ dacArea_dac_cnt_7\[4\] net57 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4925__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3774_ _3234_ _3278_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6562_ _2719_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5513_ _1694_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6493_ _2662_ _2666_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6678__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5444_ _0176_ _3084_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6142__A3 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4153__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3900__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4326_ _0177_ _3032_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4257_ _0183_ _3025_ _0372_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5653__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__A3 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4188_ _0343_ _0346_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3664__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4882__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3498__I _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5169__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6829_ _0137_ net65 dacArea_dac_cnt_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3961__I _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3407__A1 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4907__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__A2 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3490_ _3059_ net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4135__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _1347_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4111_ _0280_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5091_ _1278_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_42_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ net125 _0248_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5635__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5993_ dspArea_regP\[27\] _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6060__A2 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4944_ dspArea_regP\[15\] _1025_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4071__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4875_ _1061_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6614_ _2774_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3826_ _3317_ _3318_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6545_ dspArea_regP\[34\] _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5571__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3757_ _3264_ _3263_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3982__S _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6476_ _0213_ _3105_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3688_ dacArea_dac_cnt_3\[2\] net19 _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4126__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A1 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1611_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5174__I1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5358_ _1408_ _1543_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input43_I la_data_in[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _0213_ _3001_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5289_ _1472_ _1473_ _1474_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5626__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ net148 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3956__I _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5562__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5314__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5865__A2 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3876__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6814__A1 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5617__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3866__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4660_ _0847_ _0851_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3611_ _3118_ _3150_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _0784_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_7_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6330_ _2504_ _2505_ _2477_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3542_ _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_7_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4108__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _0226_ _3080_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3473_ _3045_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5856__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5212_ _1396_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3867__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6192_ _2312_ _2368_ _2369_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _1227_ _1229_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A2 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__A1 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _1172_ _1180_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ _0234_ net103 _0169_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6033__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__A1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _2080_ _2153_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__3398__A3 _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5792__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _0406_ _3048_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4858_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_21_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3809_ _3304_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5544__A1 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4789_ _0967_ _0970_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6528_ _2630_ _2646_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_14_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _2632_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3561__A3 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4510__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4274__A1 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6015__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _0206_ _3074_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_61_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4026__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _1844_ _1846_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _0211_ _3025_ _0734_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ _1783_ _1795_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5526__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _0192_ _3036_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4574_ _0762_ _0766_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _2268_ _2331_ _2412_ _2347_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3525_ _3087_ _3088_ net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5829__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _0197_ _3105_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3456_ dspArea_regA\[7\] _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ dspArea_regP\[29\] _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_57_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _1313_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _1182_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4008_ _0215_ _0220_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4568__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _2124_ _2138_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4740__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6245__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6860__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__A3 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3464__C1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4008__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5508__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4040__I _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4290_ _0430_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6931_ _0085_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _0016_ net65 dacArea_dac_cnt_5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5813_ _0242_ _3046_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5747__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _2936_ _2955_ _2957_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _1920_ _1921_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _1741_ _1742_ _1739_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _0816_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_2_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ _0364_ _3029_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3508_ dspArea_regA\[17\] _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4488_ _0682_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_143_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6227_ _2403_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ _3018_ net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6883__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _2164_ _2166_ _2335_ _2336_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _1294_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6089_ _2266_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5738__A1 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__I _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6466__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__I _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3790_ _3288_ _3289_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4401__A1 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5460_ _1524_ _1531_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0536_ _0539_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4704__A2 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _1411_ _1421_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4342_ _0536_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6457__A2 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4273_ _0167_ _3036_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4468__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _2190_ _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
.ends

