* NGSPICE file created from DSP48.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

.subckt DSP48 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] user_clock2 vdd vss wb_ACK wb_ADR[0] wb_ADR[10]
+ wb_ADR[11] wb_ADR[12] wb_ADR[13] wb_ADR[14] wb_ADR[15] wb_ADR[16] wb_ADR[17] wb_ADR[18]
+ wb_ADR[19] wb_ADR[1] wb_ADR[20] wb_ADR[21] wb_ADR[22] wb_ADR[23] wb_ADR[24] wb_ADR[25]
+ wb_ADR[26] wb_ADR[27] wb_ADR[28] wb_ADR[29] wb_ADR[2] wb_ADR[30] wb_ADR[31] wb_ADR[3]
+ wb_ADR[4] wb_ADR[5] wb_ADR[6] wb_ADR[7] wb_ADR[8] wb_ADR[9] wb_CYC wb_DAT_MISO[0]
+ wb_DAT_MISO[10] wb_DAT_MISO[11] wb_DAT_MISO[12] wb_DAT_MISO[13] wb_DAT_MISO[14]
+ wb_DAT_MISO[15] wb_DAT_MISO[16] wb_DAT_MISO[17] wb_DAT_MISO[18] wb_DAT_MISO[19]
+ wb_DAT_MISO[1] wb_DAT_MISO[20] wb_DAT_MISO[21] wb_DAT_MISO[22] wb_DAT_MISO[23] wb_DAT_MISO[24]
+ wb_DAT_MISO[25] wb_DAT_MISO[26] wb_DAT_MISO[27] wb_DAT_MISO[28] wb_DAT_MISO[29]
+ wb_DAT_MISO[2] wb_DAT_MISO[30] wb_DAT_MISO[31] wb_DAT_MISO[3] wb_DAT_MISO[4] wb_DAT_MISO[5]
+ wb_DAT_MISO[6] wb_DAT_MISO[7] wb_DAT_MISO[8] wb_DAT_MISO[9] wb_DAT_MOSI[0] wb_DAT_MOSI[10]
+ wb_DAT_MOSI[11] wb_DAT_MOSI[12] wb_DAT_MOSI[13] wb_DAT_MOSI[14] wb_DAT_MOSI[15]
+ wb_DAT_MOSI[16] wb_DAT_MOSI[17] wb_DAT_MOSI[18] wb_DAT_MOSI[19] wb_DAT_MOSI[1] wb_DAT_MOSI[20]
+ wb_DAT_MOSI[21] wb_DAT_MOSI[22] wb_DAT_MOSI[23] wb_DAT_MOSI[24] wb_DAT_MOSI[25]
+ wb_DAT_MOSI[26] wb_DAT_MOSI[27] wb_DAT_MOSI[28] wb_DAT_MOSI[29] wb_DAT_MOSI[2] wb_DAT_MOSI[30]
+ wb_DAT_MOSI[31] wb_DAT_MOSI[3] wb_DAT_MOSI[4] wb_DAT_MOSI[5] wb_DAT_MOSI[6] wb_DAT_MOSI[7]
+ wb_DAT_MOSI[8] wb_DAT_MOSI[9] wb_SEL wb_STB wb_WE wb_clk_i wb_rst_i
XFILLER_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6914_ _2744_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_23_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7531__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input108_I wb_DAT_MOSI[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _2579_ _2580_ _2577_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _2532_ _2535_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ _3499_ _3506_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_17_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _1567_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_13_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6145__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5658_ _1404_ _1499_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input73_I wb_ADR[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4609_ _3304_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _1344_ _1433_ _1357_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7328_ _0362_ _3461_ _3114_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6448__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7259_ _3084_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6687__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7554__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3869__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _0810_ _0765_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4622__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ _3445_ _3446_ net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4891_ _0674_ _0685_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_33_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6630_ _2310_ _2464_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A1 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3842_ _3384_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6561_ _2377_ _2379_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3773_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5512_ _1356_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ _2214_ _2216_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _0893_ _0894_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5374_ _1206_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7025__B _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ _2874_ _2870_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4325_ net123 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7044_ _1759_ _3473_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4256_ _0163_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4187_ dacArea_dac_cnt_5\[4\] net39 _3664_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_28_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3779__I _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3967__A3 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _0333_ _2493_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6366__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3719__A3 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _2591_ _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4403__I _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6118__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7577__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__I1 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5580__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4110_ dacArea_dac_cnt_3\[4\] net21 _3603_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_78_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5096__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4041_ _3548_ _3546_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6832__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4843__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6596__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5399__A2 dspArea_regA\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5992_ _1810_ _1811_ _1809_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_80_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _0730_ _0733_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7662_ net194 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6348__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4874_ dspArea_regP\[9\] _0725_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6613_ _2246_ _2250_ _2448_ _2240_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_60_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3825_ _3369_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7593_ _0113_ clknet_3_3__leaf_wb_clk_i dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6544_ _2302_ _2303_ _2308_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ dspArea_regP\[34\] _3281_ _3289_ _3308_ _3297_ dspArea_regP\[2\] _3309_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _2301_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _1185_ _1269_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6520__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4379__B _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5357_ _1113_ _1123_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0203_ _0204_ _0205_ _0206_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_59_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _1133_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input36_I la_data_in[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__I dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ dspArea_regP\[31\] _2796_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ dacArea_dac_cnt_6\[6\] net50 _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__A1 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__B _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__A2 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A3 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5002__A1 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _0444_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_31_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6750__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4978__I _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1234_ _3423_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5211_ _0264_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6191_ _2027_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_9_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5142_ _0981_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A3 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5073_ _0918_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_38_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4024_ dacArea_dac_cnt_1\[2\] net2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4292__A2 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A1 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _1813_ _1815_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5241__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ dspArea_regP\[9\] _0698_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5792__A2 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _0638_ _0641_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _3354_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7576_ _0096_ clknet_3_7__leaf_wb_clk_i dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_4788_ _0638_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6527_ _2193_ _2203_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3739_ _3293_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _2280_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5409_ _1249_ _1253_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6389_ _2128_ _2129_ _2127_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_47_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4283__A2 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6980__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7174__I _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4274__A2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5471__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__I _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5760_ _1428_ _1498_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5774__A2 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4711_ _0469_ _3329_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _1532_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7430_ _3365_ _0370_ _3247_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4642_ _0452_ _0493_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6723__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5526__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _3144_ _3146_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4573_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2148_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7292_ _3106_ _3117_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6243_ _1445_ _3403_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5829__A3 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _1895_ _1912_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ _0866_ _0867_ _0863_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_58_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _0822_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4265__A2 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4007_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3787__I _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5214__A1 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6962__A1 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _1782_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3776__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3776__B2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4909_ _0760_ _3315_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5889_ _1730_ _1664_ _1667_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5517__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7559_ _0079_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4411__I _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__I0 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4008__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__A1 dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__B2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4321__I _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4247__A2 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6930_ _2760_ _2692_ _2761_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5995__A2 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _2606_ _2607_ _2604_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5812_ _1651_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6792_ _2619_ _2622_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6795__I1 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ dspArea_regP\[17\] _1480_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ _1515_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7413_ dspArea_regP\[40\] _3234_ _0379_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4625_ dspArea_regP\[4\] _0434_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7344_ _3167_ _3168_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4183__A1 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _0414_ _0388_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4722__A3 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7460__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3930__A1 dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7275_ _0350_ _3474_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4487_ _0338_ _0351_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _0358_ _3356_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__I _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _1993_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ dspArea_regA\[12\] _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1817_ _1832_ _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4238__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _0728_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7188__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3749__A1 dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3749__B2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6163__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4174__A1 _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5910__A2 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput120 wb_DAT_MOSI[6] net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7179__A1 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4316__I _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7483__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__A1 dspArea_regP\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__I _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A2 dspArea_regA\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _1235_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4341_ _3393_ _0224_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _2802_ _2817_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4272_ dacArea_dac_cnt_7\[5\] net58 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6457__A3 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6011_ _0359_ _3340_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5665__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5968__A2 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6090__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _0361_ _3401_ _2688_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_39_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _2579_ _2580_ _2577_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_11_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3987_ dacArea_dac_cnt_0\[3\] net34 _3505_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6775_ _2566_ _2604_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_50_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6393__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _1568_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5657_ _1314_ _1500_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4608_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5588_ _1347_ _1349_ _1355_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input66_I wb_ADR[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4896__I _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7327_ _3150_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4539_ _0382_ _0393_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7258_ _3048_ _3049_ _3083_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6209_ _1936_ _2046_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7189_ _3015_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4631__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A2 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4698__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ dspArea_regP\[19\] _3429_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _0741_ _0684_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3841_ _3383_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5178__A3 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _2381_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3772_ _3322_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5511_ _1347_ _1349_ _1355_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6491_ _2214_ _2216_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7324__A1 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _0723_ _0728_ _0796_ _0878_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_8_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5373_ _1211_ _1216_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5605__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4324_ _0214_ _0216_ _0217_ _0218_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7112_ _2939_ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7025__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A1 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ _2871_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _3487_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4310__A1 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ _3662_ _3660_ _3663_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_41_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input120_I wb_DAT_MOSI[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A1 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6880__B _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _0341_ _3424_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3795__I dspArea_regA\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6758_ _0332_ _1582_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _1549_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6118__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ _2514_ _2522_ _2523_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5629__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__A3 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5801__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7521__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ dacArea_dac_cnt_1\[5\] net5 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1818_ _1827_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4942_ _0740_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7661_ net195 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4873_ _0395_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6348__A2 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ _2348_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3824_ _3368_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7592_ _0112_ clknet_3_6__leaf_wb_clk_i dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5020__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3755_ _3307_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6543_ _2285_ _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _2309_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _1099_ _1270_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6520__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5356_ _1119_ _1122_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _0193_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _1134_ _3358_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6284__A1 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ dacArea_dac_cnt_6\[6\] net50 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7026_ _3558_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I la_data_in[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ dacArea_dac_cnt_5\[0\] net35 _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5070__I dspArea_regA\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4598__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__I _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6027__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout216_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4513__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6190_ _1838_ _2028_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _0896_ _0982_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _0919_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4816__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4023_ _3516_ _3534_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6018__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _1813_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5241__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4925_ _0774_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_80_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7567__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4856_ _0686_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3807_ _3353_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7575_ _0095_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4787_ _0569_ _0639_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3738_ _3292_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5065__I _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6457_ _2285_ _2290_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_69_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5552__I0 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _1151_ _1153_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6388_ _2190_ _2222_ _2225_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5339_ _1096_ _1097_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6257__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _2823_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4409__I _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4283__A3 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_18_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6980__A2 dspArea_regA\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5299__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4319__I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__A2 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4054__I _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _0564_ _3322_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ _1533_ _3317_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4641_ _0337_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6723__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4734__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7360_ _3175_ _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4572_ _0428_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6311_ _2055_ _2067_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7291_ _3108_ _3116_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_6_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6242_ _1443_ _3395_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _1907_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _0934_ _0970_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_5055_ _0902_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_57_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ _3490_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _1795_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4973__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _0615_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5888_ _1573_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input96_I wb_ADR[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4839_ _0687_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6714__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _0078_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _2166_ _2344_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ _0009_ net213 dacArea_dac_cnt_4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6478__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6619__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6650__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__I1 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3978__I _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3767__A2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7130__A2 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6641__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3888__I _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _2676_ _2679_ _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_23_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _1652_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6791_ _2246_ _2250_ _2623_ _2624_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ _1583_ _1585_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5673_ _1516_ _1427_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7412_ _3225_ _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4624_ _0475_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7343_ _3142_ _3143_ _3166_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5380__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _0386_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7274_ _0343_ _3482_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _0350_ net103 _0344_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6225_ _2062_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5343__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _1994_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _0570_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ _1835_ _1927_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_57_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6632__A1 dspArea_regB\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _0883_ _0884_ _0886_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I la_data_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7188__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6989_ _2714_ _2716_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_80_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3749__A2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I dspArea_regB\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5371__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput110 wb_DAT_MOSI[1] net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_1_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput121 wb_DAT_MOSI[7] net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6623__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6926__A2 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4332__I _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7351__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ net103 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4271_ _0164_ _0176_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5163__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input3_I la_data_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7311__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6912_ _0356_ _3410_ _2686_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_82_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _2675_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4928__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _2606_ _2607_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3986_ dacArea_dac_cnt_0\[2\] net23 _3504_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5725_ _0296_ _1059_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _1383_ _1386_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4156__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _0282_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5587_ _1326_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7326_ _1406_ _3469_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_2_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4538_ _0364_ _0397_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input59_I la_data_in[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7257_ _3048_ _3049_ _3083_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_46_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _0335_ net101 _0316_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _2024_ _2025_ _2021_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7188_ _1845_ _3451_ _2949_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6139_ _1342_ _3399_ _1890_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4417__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5344__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4083__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ dspArea_regA\[12\] _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5158__I _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _1347_ _1349_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_34_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6490_ _2209_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7324__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5441_ _1275_ _1282_ _1283_ _1284_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5372_ _1217_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _1333_ _3473_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _0193_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _0327_ _3467_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4254_ _3692_ _0162_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4185_ dacArea_dac_cnt_5\[3\] net38 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input113_I wb_DAT_MOSI[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__A2 dspArea_regA\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _1305_ _3416_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _0341_ _1478_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3969_ _3490_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _1550_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6688_ _1775_ _3465_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7315__A2 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5639_ _1366_ _1370_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__I dspArea_regA\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _3133_ _3134_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_output165_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6826__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7473__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7003__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A3 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7306__A2 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4540__A2 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout196_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _0987_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _0789_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3896__I _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ net196 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4872_ _0723_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6348__A3 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6611_ _2444_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5556__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3823_ _3367_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7591_ _0111_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6542_ _2290_ _2293_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3754_ _3306_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _2302_ _2303_ _2308_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5424_ _1166_ _1169_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5355_ _1186_ _1189_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__5552__S _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4306_ _3326_ _0201_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7496__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5286_ dspArea_regB\[5\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7025_ _2784_ _2454_ _2854_ _2855_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6284__A2 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4237_ _3692_ _3704_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5351__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4168_ dacArea_dac_cnt_5\[0\] net35 _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4099_ dacArea_dac_cnt_3\[2\] net19 _3594_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_55_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4598__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6809_ _2640_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4430__I _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4522__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__I _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6027__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6092__I _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__I _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4340__I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout209_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4513__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7651__I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5140_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_9_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5071_ _0313_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_57_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ dacArea_dac_cnt_1\[2\] net2 _3533_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4816__A3 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7215__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _1626_ _1713_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_52_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4924_ dspArea_regP\[10\] _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _0704_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_18_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _3352_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7574_ _0094_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4786_ _0574_ _0576_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6525_ _2269_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3737_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4752__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _2291_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5407_ dspArea_regP\[14\] _1152_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5701__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__I1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _2223_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5338_ _1092_ _1098_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input41_I la_data_in[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6257__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _1116_ dspArea_regA\[6\] _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7008_ _2827_ _2838_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_47_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__I _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7511__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__B _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5940__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7445__A1 _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _0451_ _0494_ _0496_ _0261_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6723__A3 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4571_ _0292_ _3292_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5931__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6310_ _2058_ _2066_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7290_ _3114_ _3115_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6487__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _0325_ _3390_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6172_ _1910_ _1915_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_44_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7436__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _0971_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5054_ _0809_ _0903_ _0902_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5998__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ _3516_ _3520_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7534__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5956_ _1689_ _1796_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _0757_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4973__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5887_ _1564_ _1574_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4838_ _0688_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6175__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input89_I wb_ADR[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7557_ _0077_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5076__I dspArea_regB\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _2226_ _2229_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7488_ _0008_ net210 dacArea_dac_cnt_4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6478__A2 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6439_ _2182_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__A2 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7427__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6650__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4661__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4155__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7557__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6641__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5810_ _1109_ dspArea_regA\[8\] _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6790_ _2441_ _2542_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6944__A3 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ dspArea_regP\[18\] _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5672_ _1409_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7411_ _3229_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ dspArea_regP\[5\] _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5904__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7342_ _3142_ _3143_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_4554_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5380__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7273_ dspArea_regP\[35\] _3057_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4485_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6224_ _2059_ _2060_ _2061_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _0276_ dspArea_regA\[20\] _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1838_ _1923_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _0885_ _0721_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6632__A2 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6988_ _2798_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_40_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _1779_ _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6404__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6148__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5371__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6320__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput100 wb_DAT_MOSI[10] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput111 wb_DAT_MOSI[20] net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput122 wb_DAT_MOSI[8] net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4882__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6623__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4270_ dacArea_dac_cnt_7\[5\] net58 _0175_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6275__I _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4625__A1 dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6911_ _2737_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _2652_ _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_36_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ _2501_ _2531_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3985_ _3501_ _3503_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5724_ _0507_ _0959_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _1383_ _1386_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4606_ _0460_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5586_ _1331_ _1335_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7325_ _3148_ _0355_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4537_ dspArea_regP\[2\] _0394_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5354__I _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7256_ _3076_ _3079_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6302__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6207_ _2024_ _2025_ _2021_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7187_ _0343_ _3468_ _2866_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4399_ _0262_ _0275_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6138_ _1225_ _1884_ _1776_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6605__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6069_ _1791_ _1793_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__A2 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A2 _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__I _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4343__I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3770_ dspArea_regA\[4\] _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7654__I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5440_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6532__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _0326_ _0433_ _1118_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7110_ _1759_ _3479_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4322_ _3356_ _0212_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7041_ _2869_ _2870_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4253_ dacArea_dac_cnt_7\[2\] net54 _0161_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4846__A1 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4184_ dacArea_dac_cnt_5\[3\] net38 _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4518__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input106_I wb_DAT_MOSI[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _2656_ _2657_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5023__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ net126 _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6756_ _1013_ _3407_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_32_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1022_ _1038_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6687_ dspArea_regB\[7\] _2108_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3899_ _3435_ _3418_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5638_ dspArea_regP\[16\] _1369_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input71_I wb_ADR[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7308_ _3132_ _3093_ _3098_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_144_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6826__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ _2948_ _3052_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_63_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4837__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4428__I dspArea_regB\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6643__I _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7003__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4338__I _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7649__I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _0669_ _0790_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4871_ _0659_ _0661_ _0722_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5169__I dspArea_regB\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _2235_ _2238_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_60_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3822_ _3366_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7590_ _0110_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6541_ _2290_ _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3753_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6472_ _2302_ _2303_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _1166_ _1169_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _0189_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6808__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5285_ _0507_ _1045_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4819__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7024_ _3490_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4236_ dacArea_dac_cnt_6\[6\] net50 _3703_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4295__A2 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4167_ _3645_ _3649_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4098_ _3593_ _3592_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__A3 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _1775_ _2319_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6739_ _0297_ _2210_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3730__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7590__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7224__A2 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4038__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6735__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4621__I _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5070_ dspArea_regA\[4\] _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4277__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__I _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ _3532_ _3531_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7215__A2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4029__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6974__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _1709_ _1712_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_64_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _0264_ _3366_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _0630_ _0705_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ dspArea_regA\[8\] _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7573_ _0093_ clknet_3_7__leaf_wb_clk_i dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4785_ _0574_ _0576_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4201__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4531__I _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _1405_ _3371_ _2270_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3736_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7463__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3960__A1 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6455_ _1970_ _3398_ _2181_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5406_ _1250_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6386_ _2106_ _2126_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5701__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5337_ _1089_ _1182_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5268_ dspArea_regB\[8\] _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6257__A3 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4268__A2 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I la_data_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ dacArea_dac_cnt_6\[2\] net46 _3689_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7007_ _2830_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _1043_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__I _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6717__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4441__I _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7142__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4259__A2 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7381__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__I _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout221_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4570_ _0409_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7662__I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _2075_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6171_ _1991_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _0845_ _0862_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7436__A2 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5053_ _0813_ _0826_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5998__A2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7103__S _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4004_ dacArea_dac_cnt_0\[6\] net61 _3519_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _1693_ _1695_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _0678_ _3331_ _0691_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5886_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _0277_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7372__A1 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7556_ _0076_ clknet_3_6__leaf_wb_clk_i dspArea_regB\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ dspArea_regB\[4\] _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6507_ _2226_ _2229_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3719_ net77 net66 _3272_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7487_ _0007_ net212 dacArea_dac_cnt_4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4699_ dspArea_regB\[5\] _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6438_ _2185_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _0468_ dspArea_regA\[22\] _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_1_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A2 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4436__I _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A1 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4346__I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__A2 dspArea_regA\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7657__I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5601__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ _0476_ dspArea_regA\[18\] _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5671_ _1412_ _1426_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7410_ dspArea_regP\[40\] _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4622_ _0477_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5904__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7341_ _3161_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4553_ _0406_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5380__A3 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _3094_ _3095_ _3097_ _3085_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4484_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5668__A1 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _2059_ _2060_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7501__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _1244_ dspArea_regA\[19\] _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ dspArea_regA\[11\] _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _1741_ _1924_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_58_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _0885_ _0721_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_2_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5840__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4256__I _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6987_ _2802_ _2817_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6396__A2 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5938_ _1771_ _1772_ _1778_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6404__C _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A2 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _1537_ _1710_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7539_ _0059_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6320__A2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_DAT_MOSI[11] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput112 wb_DAT_MOSI[21] net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput123 wb_DAT_MOSI[9] net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4882__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6084__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A1 dspArea_regB\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A2 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4322__A1 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6910_ _2740_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6841_ _2655_ _2658_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_1_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _2605_ _2530_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ dacArea_dac_cnt_0\[2\] net23 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5723_ _0551_ _3376_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5654_ _1428_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4605_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_15_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6550__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _1331_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7324_ _3052_ _3145_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_7_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4536_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7255_ _3080_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4313__A1 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _1831_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7186_ _3013_ _2955_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4398_ _0274_ net110 _0269_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _1975_ _1976_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6068_ _1791_ _1793_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ _0786_ _0787_ _0785_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__A2 dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6844__A3 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4791__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6532__A2 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4543__A1 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0321_ _3337_ _1023_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4321_ _0215_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7670__I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _0160_ _0159_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7040_ _0314_ _2319_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4846__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ _3639_ _3661_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5190__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6048__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6824_ _2571_ _2575_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _2587_ _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3967_ net124 net98 _3489_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_50_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _0319_ _3358_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4782__A1 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _2518_ _2519_ _2520_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3898_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ _1479_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5568_ _0915_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input64_I la_data_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7307_ _3093_ _3098_ _3132_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4519_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5499_ _0284_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7238_ _3064_ _3005_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_78_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _0334_ _3474_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6762__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4773__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7423__C _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4828__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__I _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6450__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4354__I _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ _0659_ _0661_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ dspArea_regA\[10\] _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7665__I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4764__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _2293_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3752_ _3304_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6471_ _2304_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6505__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _1202_ _1265_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5353_ _1196_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_47_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5913__I _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ net118 _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5284_ _0306_ _3345_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7023_ _1831_ _2852_ _2853_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4235_ dacArea_dac_cnt_6\[5\] net49 _3702_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4166_ net195 net33 _3648_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_67_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ dacArea_dac_cnt_3\[1\] net18 _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6807_ _0839_ _3472_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4999_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4755__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _0305_ _3456_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _2502_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4507__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5180__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3730__A2 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6432__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A2 _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__A2 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A3 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5171__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ dacArea_dac_cnt_1\[1\] net64 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6671__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _1725_ _1809_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6974__A2 _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ _0272_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4853_ _0635_ _0637_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_18_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3804_ _3280_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7572_ _0092_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4784_ _0630_ _0635_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _2356_ _2358_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3735_ dspArea_regA\[0\] _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3960__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _1968_ _3415_ _2082_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7151__A2 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ dspArea_regP\[15\] _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _2122_ _2125_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5336_ _1170_ _1172_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _0735_ dspArea_regA\[5\] _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7006_ _2835_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5465__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6662__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4218_ _3686_ _3688_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5198_ _1044_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input27_I la_data_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4149_ _3623_ _3634_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6965__A2 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6717__A2 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5776__I0 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7142__A2 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4900__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5208__A2 _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6708__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7381__A2 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4195__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6892__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _2005_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5121_ _0857_ _0861_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6644__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _0813_ _0826_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4003_ dacArea_dac_cnt_0\[5\] net56 _3518_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4958__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _1693_ _1695_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _0627_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5885_ _1639_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4836_ _3343_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7555_ _0075_ clknet_3_6__leaf_wb_clk_i dspArea_regB\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5383__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _0610_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7580__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6506_ _2274_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3718_ net97 net96 net68 net67 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7486_ _0006_ net212 dacArea_dac_cnt_4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _0551_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5135__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6437_ _2261_ _2273_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6883__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6368_ _0282_ _2110_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5319_ _1071_ _1072_ _1070_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6299_ _2136_ _2137_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6635__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7060__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__A1 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6626__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7453__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__A2 dspArea_regA\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _3498_ _1399_ _1514_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4621_ _3328_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5365__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4412__I0 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5904__A3 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _3162_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4552_ _0407_ _0408_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7271_ _3088_ _3096_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4483_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6222_ _1636_ _3362_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6153_ _0289_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _1805_ _1808_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4479__I0 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6093__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _0717_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7042__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6986_ _2803_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_53_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5937_ _1771_ _1772_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5868_ _1598_ _1601_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A3 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input94_I wb_ADR[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ _0556_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5356__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _1640_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7538_ _0058_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7469_ _0143_ net205 dacArea_dac_cnt_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6856__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__A3 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput102 wb_DAT_MOSI[12] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput113 wb_DAT_MOSI[22] net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput124 wb_STB net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7476__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5831__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5898__A2 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6847__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7668__I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _2663_ _2672_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2527_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3983_ _3499_ _3502_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1348_ _1346_ _1475_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_15_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7327__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5653_ _1494_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_30_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4604_ _3299_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5584_ _1335_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _0355_ _3475_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4535_ _0369_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7254_ _3012_ _3022_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4466_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7499__CLK net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6205_ dspArea_regP\[23\] _1085_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5510__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ _2951_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4397_ _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _1953_ _1955_ _1974_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__A1 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6067_ _1787_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _0827_ _0863_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6482__I dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6969_ _2731_ _2733_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_10_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__I _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__A1 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5804__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5740__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _0188_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4251_ dacArea_dac_cnt_7\[1\] net53 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4182_ dacArea_dac_cnt_5\[3\] net38 _3660_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_67_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I la_data_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7245__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6048__A2 _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__B _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _2506_ _2574_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__A2 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6754_ _2517_ _2525_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3966_ _3488_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5705_ _1019_ _0695_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6685_ _0279_ _3479_ _2404_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4782__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _3433_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5636_ dspArea_regP\[17\] _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5731__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _1411_ _1336_ _1339_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7306_ _3127_ _3131_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4518_ _0369_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _1341_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input57_I la_data_in[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _3001_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6477__I dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6287__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ dspArea_regB\[9\] _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _0342_ _3467_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6039__A2 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _1437_ _1038_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7099_ _2242_ _2245_ _2926_ _2927_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5798__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7514__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4773__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__I _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6278__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3804__I _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4289__A1 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7227__A1 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6450__A2 _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ dspArea_regP\[42\] _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3751_ dspArea_regA\[2\] _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4764__A2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _2305_ _2306_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5421_ _1126_ _1266_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5713__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5352_ _1198_ _0390_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ _0199_ _0190_ _0202_ _0194_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5283_ _0291_ _3360_ _1054_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _2786_ _2788_ _2851_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4234_ _3701_ _3699_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_4_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4165_ _3646_ _3643_ _3647_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7537__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4096_ _3559_ _3591_ _3592_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input111_I wb_DAT_MOSI[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _1886_ _3466_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4204__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ _0846_ _0847_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _3479_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6737_ _2522_ _2568_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4755__A2 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5952__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6668_ _0624_ _2210_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5619_ _1234_ _3375_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6599_ _2274_ _2342_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6432__A2 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A3 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6196__A1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__I dspArea_regB\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7448__A1 _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout194_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6423__A2 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _1810_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _3359_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _0635_ _0637_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6187__A1 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3803_ _3350_ net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7571_ _0091_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_18_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4737__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5196__I dspArea_regA\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _0571_ _0573_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5934__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _2357_ _2273_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3734_ _3288_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _2286_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5404_ _0697_ _3404_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6384_ _2204_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7439__A1 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5335_ _1170_ _1172_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5266_ _1018_ _3321_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6111__A1 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7005_ _1424_ _3417_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4217_ dacArea_dac_cnt_6\[2\] net46 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6662__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5197_ _0295_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ dacArea_dac_cnt_4\[4\] net30 _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_55_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4079_ dacArea_dac_cnt_2\[5\] net14 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6965__A3 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__I _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__I1 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7142__A3 _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4900__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6102__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__C1 _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6405__A2 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout207_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6892__A2 _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _0948_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5051_ _0808_ _0899_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4655__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4002_ _3517_ _3513_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_38_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ _1787_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4904_ _0564_ _3344_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5884_ _1406_ _3326_ _1640_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5907__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _0464_ _3336_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7554_ _0074_ clknet_3_6__leaf_wb_clk_i dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6580__A1 dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _0613_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5383__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3717_ net70 net69 net72 net71 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_6505_ _2338_ _2341_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7485_ _0005_ net210 dacArea_dac_cnt_4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4697_ dspArea_regA\[0\] _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6436_ _2264_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6332__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6367_ _0561_ _3448_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4894__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5318_ _1126_ _1162_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6298_ _1951_ _2020_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__A2 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _0355_ _0391_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7521__D _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3902__I dspArea_regA\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4646__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5071__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6571__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6626__A2 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4908__I _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3812__I dspArea_regA\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__C1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5062__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5365__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4412__I1 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4551_ _0392_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_7270_ _3084_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4482_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6221_ _1634_ _3362_ _1961_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _3431_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0950_ _0951_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6617__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _1805_ _1808_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4479__I1 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _0660_ _0652_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7042__A2 _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _2808_ _2813_ _2815_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_81_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5936_ _1773_ _1777_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4800__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _1598_ _1601_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6553__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _0301_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5356__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _1198_ _3326_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input87_I wb_ADR[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7537_ _0057_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4749_ _0601_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7468_ _0142_ net203 dacArea_dac_cnt_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6856__A2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6419_ _2150_ _2234_ _2255_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7399_ _3098_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_1_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput103 wb_DAT_MOSI[13] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput114 wb_DAT_MOSI[23] net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput125 wb_WE net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6544__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3807__I _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4858__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4638__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__A3 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7570__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5469__I _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3982_ dacArea_dac_cnt_0\[2\] net23 _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6770_ _2577_ _2581_ _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5721_ _1345_ _3408_ _1362_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _1340_ _1495_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _0290_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5583_ _1409_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4534_ _0382_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7322_ _3144_ _3146_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _3014_ _3021_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4465_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6204_ _1932_ _2043_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7184_ _3010_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4396_ _0272_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5510__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _1953_ _1955_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _1900_ _1904_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6066__A3 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _0866_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ _2726_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ _0748_ _3361_ _1659_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6899_ _2727_ _2730_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5501__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4458__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7593__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4921__I _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7190__A1 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5740__A2 dspArea_regA\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _3681_ _0158_ _0159_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6296__A3 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ dacArea_dac_cnt_5\[2\] net37 _3659_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_68_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7245__A2 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6822_ _2594_ _2653_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_1_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6756__A1 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3965_ _3487_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4231__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _1544_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6684_ _2404_ _2419_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3896_ _3432_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5635_ _0697_ _3422_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _1240_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_3_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7305_ _3128_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4517_ _0373_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_2_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4479__S _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5497_ _1342_ _3354_ _1237_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7236_ _3061_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _0311_ _0317_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4298__A2 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7167_ _1845_ _3460_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4379_ _0257_ _0250_ _0258_ _0252_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _0346_ _3359_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6039__A3 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2923_ _2926_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _1888_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_73_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6995__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5798__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7172__A1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4289__A2 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5486__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4916__I dspArea_regB\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7489__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__I dspArea_regB\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3750_ _3303_ net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _1163_ _1164_ _1162_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3724__A1 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4302_ _3317_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5282_ _0547_ _0956_ _0952_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4233_ dacArea_dac_cnt_6\[5\] net49 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7021_ _2786_ _2788_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_4_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ dacArea_dac_cnt_4\[6\] net32 _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4095_ _3589_ _3590_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6977__A1 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6729__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input104_I wb_DAT_MOSI[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6805_ dspArea_regP\[29\] _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4997_ _0279_ _3360_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _2409_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3948_ _3478_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5952__A2 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3963__A1 dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _0284_ _3479_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3879_ _3310_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5618_ _0615_ _3368_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6901__A1 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _2338_ _2341_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5549_ _1092_ _1098_ _1393_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__I _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _2856_ _3046_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_28_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4691__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4471__I _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A1 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7145__A1 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__I _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A1 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _0756_ _0770_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _0693_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_60_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3802_ dspArea_regP\[39\] _3320_ _3342_ _3348_ _3349_ dspArea_regP\[7\] _3350_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7570_ _0090_ clknet_3_3__leaf_wb_clk_i dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4782_ dspArea_regP\[7\] _0572_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5934__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3945__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _2261_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3733_ _3287_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6452_ _2287_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5403_ _0694_ _3397_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6383_ _2217_ _2220_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7504__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5334_ dspArea_regP\[15\] _0799_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_47_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5265_ _1108_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7004_ _2833_ _2834_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4216_ _3666_ _3687_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ dspArea_regA\[8\] _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4147_ _3631_ _3629_ _3632_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4078_ _3570_ _3578_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5622__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7519__D _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4291__I _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6719_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6102__A2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__I _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__B1 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3872__C2 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5613__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7218__S _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7527__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6341__A2 _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4352__A1 _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5050_ _0869_ _0872_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_46_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ dacArea_dac_cnt_0\[5\] net56 _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4655__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5604__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _1791_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ _0753_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ _1722_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _0677_ _0521_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5907__A2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7553_ _0073_ clknet_3_6__leaf_wb_clk_i dspArea_regB\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4765_ _0616_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6580__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5383__A3 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _2190_ _2339_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4591__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3716_ _3266_ _3270_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7484_ _0004_ net210 dacArea_dac_cnt_4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4696_ _0305_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_14_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _2270_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6366_ _2193_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_88_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4894__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5317_ _1163_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _2016_ _2019_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_25_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5248_ _1094_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input32_I la_data_in[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__I _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4646__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__A1 dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _1026_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6399__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6020__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3909__A1 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6571__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7265__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__C _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__I0 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5834__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__B1 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3845__C2 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4550_ _0285_ _3300_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ dspArea_regB\[13\] _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6220_ _1632_ _3378_ _1864_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _1980_ _1990_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5102_ _0278_ _3367_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _1855_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0597_ _0656_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6984_ _2727_ _2730_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5935_ _1774_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5866_ _1644_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _3313_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5797_ _1638_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6553__A2 dspArea_regA\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7536_ _0056_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4748_ _0315_ _3291_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7467_ _0141_ net204 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4679_ _0484_ _0487_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6418_ _2230_ _2233_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7398_ _3132_ _3169_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _2172_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__C _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput104 wb_DAT_MOSI[14] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput115 wb_DAT_MOSI[24] net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput126 wb_rst_i net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__C2 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__I _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6792__A2 _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5776__S _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6544__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3818__C2 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5283__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6232__A1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3981_ _3500_ _3497_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _1562_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5651_ _1380_ _1381_ _1379_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4602_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5582_ _1412_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_7_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7321_ dspArea_regP\[37\] _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4533_ _0389_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_8_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _3077_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4464_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6203_ dspArea_regP\[22\] _2042_ _1619_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7183_ _2975_ _2976_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4395_ _0271_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _1957_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _1788_ _1790_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6471__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5016_ _0767_ _0784_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_39_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__B _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5026__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2793_ _2797_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_59_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5918_ _1759_ _3377_ _1551_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6898_ _2728_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ dspArea_regP\[19\] _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3908__I _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7527__D _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7519_ _0039_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4474__I _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6214__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6765__A2 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7190__A2 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _3656_ _3658_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_79_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__I _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6205__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _2599_ _2600_ _2598_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6756__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6752_ _2521_ _2524_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3964_ net126 _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _1545_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _2418_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6508__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3895_ _3431_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ _0694_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3990__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ _1228_ _1241_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7304_ _3129_ _3082_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4516_ _0375_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5496_ _0615_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7235_ _3019_ _3020_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4447_ _0315_ net122 _0316_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5495__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ dspArea_regP\[33\] _2956_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ _3475_ _0189_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6117_ _1882_ _1956_ _1893_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _2619_ _2622_ _2922_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_59_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6444__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _1352_ _3413_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6995__A2 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7560__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4930__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6617__C _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6986__A2 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6738__A2 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4749__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3972__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5174__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5713__A3 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3724__A2 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ dspArea_regB\[15\] _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _0200_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6795__S _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _1127_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _2850_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _3692_ _3700_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ dacArea_dac_cnt_4\[6\] net32 _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4094_ _3589_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_67_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__A2 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6804_ dspArea_regP\[28\] _2505_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_63_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__I _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ _0561_ _3345_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6735_ _0604_ _2314_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3947_ dspArea_regA\[24\] _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7583__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3963__A2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6666_ _2499_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3878_ _3416_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5165__A1 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _0678_ _1229_ _1363_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6597_ _2375_ _2429_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4507__A4 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6901__A2 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3715__A2 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ _1269_ _1272_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input62_I la_data_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5479_ _1322_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ dspArea_regP\[34\] _3045_ _2628_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7149_ _2970_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4979__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5640__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7145__A2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__A1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3831__I _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__A1 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7456__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3890__A1 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _0700_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3801_ _3296_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4198__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _0632_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ _2264_ _2272_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3732_ _3285_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6451_ _1445_ dspArea_regA\[17\] _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6895__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5698__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6382_ _2114_ _2218_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5333_ _0451_ _1179_ _1180_ _1087_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__4370__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__A1 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5264_ _1093_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7003_ _1419_ _3427_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4215_ dacArea_dac_cnt_6\[2\] net46 _3686_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4122__A2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3741__I _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _0300_ _0689_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5870__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4146_ dacArea_dac_cnt_4\[3\] net29 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ dacArea_dac_cnt_2\[5\] net14 _3577_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_37_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7375__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ _0829_ _3331_ _0682_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6718_ _2472_ _2551_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7127__A2 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6649_ _1011_ _3396_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3916__I _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7479__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5861__A2 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A1 dspArea_regP\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3872__B2 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5613__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4482__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7118__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3826__I _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4352__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6629__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4000_ _3515_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6801__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _1690_ _1692_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4902_ _0309_ _3306_ _0683_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_52_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5882_ _1723_ _1643_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7357__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _0674_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_60_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6821__B _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7552_ _0072_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4764_ _0605_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6503_ _2223_ _2224_ _2222_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3715_ _3267_ _3268_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7483_ _0003_ net206 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3736__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _0548_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6112__I _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _0359_ _3371_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6365_ _2201_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5316_ _1050_ _1069_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2068_ _2131_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5247_ _0350_ _0390_ _1016_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A2 dspArea_regA\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5178_ _0928_ _0466_ _0922_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA_input25_I la_data_in[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _3587_ _3617_ _3618_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_21_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4582__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7284__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__I1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_260 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_48_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__A1 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3845__B2 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7036__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6011__A2 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5770__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout212_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _0338_ _0345_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _1988_ _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7275__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ _0768_ _0695_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4387__I _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1919_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5032_ _0337_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7027__A1 dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _0315_ _3467_ _2728_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_53_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5934_ _1775_ _3405_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4261__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ _1704_ _1707_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7604_ _0124_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _0666_ _0667_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5796_ _1633_ _1635_ _1637_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7535_ _0055_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4564__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _0599_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7466_ _0140_ net204 dacArea_dac_cnt_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4678_ _0512_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6417_ dspArea_regP\[25\] _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7397_ _3193_ _3215_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6348_ _2177_ _2182_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_27_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__A2 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput105 wb_DAT_MOSI[15] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6279_ _2115_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xinput116 wb_DAT_MOSI[2] net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3827__B2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7517__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4760__I dspArea_regB\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A3 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5504__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4000__I _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3818__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3818__B2 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ dacArea_dac_cnt_0\[1\] net12 _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5650_ _1380_ _1381_ _1379_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_31_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ _0456_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_15_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5581_ _1423_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5743__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7320_ _2893_ _3482_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _0280_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ _3008_ _3023_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6299__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4463_ dspArea_regB\[11\] _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6202_ _2031_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _3009_ _2974_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4394_ dspArea_regB\[1\] _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _1962_ _1967_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ dspArea_regP\[20\] _1789_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _0780_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7420__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ dspArea_regP\[31\] _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _0737_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4785__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ _1755_ _2314_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5848_ _1367_ dspArea_regA\[19\] _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input92_I wb_ADR[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5734__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _1603_ _1604_ _1602_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_5_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7518_ _0038_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7449_ dspArea_regP\[47\] _3263_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7543__D _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__I _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7239__A1 _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__A2 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A1 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3834__I _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _2599_ _2600_ _2598_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4216__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3963_ dspArea_regP\[31\] _3420_ net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6751_ _2582_ _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5496__I _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _0331_ _3343_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6682_ _2515_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3894_ dspArea_regA\[18\] _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5633_ _3414_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5716__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _1309_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_8_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7303_ _3076_ _3079_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4515_ _0274_ _3293_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ _1033_ _3369_ _1135_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_7234_ _3060_ _3018_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4446_ _0268_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6141__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _2934_ _2454_ _2993_ _2855_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5495__A3 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4377_ net114 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6116_ _1883_ _1885_ _1891_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7096_ _2849_ _2924_ _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4575__I _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__A2 _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6047_ _0604_ _3405_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4207__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6949_ _2777_ _2780_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5707__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7172__A3 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4694__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__I _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4749__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6371__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__A2 dspArea_regA\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _0187_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6123__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ _1043_ _1047_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4231_ dacArea_dac_cnt_6\[5\] net49 _3699_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4685__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4162_ _3491_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4395__I _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ dacArea_dac_cnt_3\[1\] net18 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_67_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _2634_ _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5937__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__I _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4995_ _0283_ _3353_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _2514_ _2523_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3946_ _3476_ _3477_ net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ _3415_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6665_ _2479_ _2481_ _2498_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_17_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _0675_ _3399_ _1246_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5165__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _2298_ _2430_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3715__A3 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5547_ _1269_ _1272_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6114__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5478_ _1323_ _3328_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input55_I la_data_in[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7217_ _3037_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4429_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4676__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7148_ _2975_ _2976_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_24_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7079_ _2827_ _2838_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_46_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4979__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4600__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6353__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5104__I _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5919__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3800_ _3347_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4780_ dspArea_regP\[8\] _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3731_ net92 _3277_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6450_ _1443_ _3413_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ _1243_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6895__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _2118_ _2120_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5332_ dspArea_regP\[14\] _0495_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__A2 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ _1110_ _3313_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4214_ _3685_ _3684_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7002_ _2831_ _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5442__C _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5194_ _0305_ _0769_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4145_ dacArea_dac_cnt_4\[3\] net29 _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _3575_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7550__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6583__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6717_ _1519_ _3387_ _2473_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3929_ _3411_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5138__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6648_ _2402_ _2482_ _2413_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6335__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _2402_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4897__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3932__I dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5613__A3 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3842__I _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout192_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__S _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6801__A2 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A3 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5950_ dspArea_regP\[19\] _1691_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0303_ _3325_ _0617_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_52_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _1628_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4832_ _0680_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5368__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7551_ _0071_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _0554_ _3313_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_53_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4040__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _2223_ _2224_ _2222_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3714_ net87 net86 net90 net89 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7482_ _0002_ net215 dacArea_dac_cnt_3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4694_ _0291_ _3305_ _0518_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _2268_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6364_ _2194_ _2195_ _2200_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5315_ _1065_ _1068_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3752__I _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6295_ _1977_ _2132_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ _0914_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_25_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _0321_ _0433_ _0817_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ dacArea_dac_cnt_4\[0\] net26 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7045__A2 _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input18_I la_data_in[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ dacArea_dac_cnt_2\[1\] net9 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6556__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6308__A1 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7596__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7284__A2 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_250 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__5295__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_261 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_48_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7036__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4270__A2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A1 dspArea_regB\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4022__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout205_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ _0564_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7275__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _1767_ _1804_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5031_ _3681_ _0800_ _0881_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_6_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7027__A2 _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5499__I _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2809_ _2812_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_81_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _1134_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6538__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5864_ _1561_ _1705_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _0123_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7469__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ _0323_ _0391_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5795_ _1633_ _1635_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7534_ _0054_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _0509_ _0559_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7465_ _0139_ net206 dacArea_dac_cnt_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4677_ _0529_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ _1932_ _2253_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6710__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _3199_ _0423_ _3218_ _3521_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _2183_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6278_ dspArea_regP\[23\] _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xinput106 wb_DAT_MOSI[16] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput117 wb_DAT_MOSI[3] net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _1074_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6777__A1 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4004__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5752__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5504__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__A2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6768__A1 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _0298_ _3290_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5580_ _1424_ _3308_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_54_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4531_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_8_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7250_ _2994_ _3007_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4462_ _0311_ _0329_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6201_ _2038_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7181_ _2973_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4393_ _0262_ _0270_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _1969_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _1901_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_58_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _0782_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_6_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _2794_ _2795_ _2640_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_53_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _1753_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6896_ _0736_ _2110_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _0271_ _3432_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5734__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5778_ _1603_ _1604_ _1602_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input85_I wb_ADR[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7517_ _0037_ clknet_3_1__leaf_wb_clk_i dspArea_regA\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4729_ _0512_ _0582_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_5_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7448_ _0154_ _3262_ _3263_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7379_ _3133_ _3194_ _3193_ _3201_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__4101__I _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7239__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4170__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__I dspArea_regA\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5670__A1 _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7175__A1 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5725__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4161__A1 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3850__I _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5413__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _2487_ _2583_ _2582_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_63_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3962_ dspArea_regP\[30\] _3420_ net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _0340_ _3335_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7166__A1 dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6681_ _0760_ _3442_ _2410_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3893_ _3428_ _3430_ net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5632_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6913__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5563_ _1407_ _3302_ _1310_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7507__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7302_ _3076_ _3079_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4514_ dspArea_regP\[1\] _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5494_ _1338_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7233_ _3017_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4445_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6141__A2 _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7164_ _1831_ _2991_ _2992_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4376_ _0255_ _0250_ _0256_ _0252_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_8_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _1866_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _2786_ _2848_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3760__I dspArea_regA\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _1886_ _3398_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2619_ _2622_ _2625_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_53_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5955__A2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6879_ _0298_ _3480_ _2640_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5707__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__I _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5946__A2 _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3957__A1 dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4006__I _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7320__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6123__A2 _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ _3697_ _3698_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4161_ _3639_ _3644_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4092_ _3587_ _3588_ _3589_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_83_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5634__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _2553_ _2565_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5937__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4994_ _0832_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6733_ dspArea_regP\[28\] _2505_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3945_ dspArea_regP\[23\] _3463_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _2479_ _2481_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3876_ _3414_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _1458_ _1459_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3755__I _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _2335_ _2336_ _2332_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5546_ _1296_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7311__A1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ dspArea_regB\[11\] _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6114__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4125__A1 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _3038_ _3040_ _3043_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4428_ dspArea_regB\[6\] _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5873__A1 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input48_I la_data_in[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7147_ _1297_ _3435_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4359_ net108 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7078_ _2830_ _2837_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _1868_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5210__I _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A2 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4739__I0 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__A2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4364__A1 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4116__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__I _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5616__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A2 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6216__I _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _3271_ _3274_ _3284_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4355__A1 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _1245_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6380_ _2118_ _2120_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5331_ _1174_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6886__I _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6647__A3 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5262_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7001_ _0349_ _3426_ _2725_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5855__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ dacArea_dac_cnt_6\[1\] net44 _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5193_ _0951_ _1037_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__C _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4144_ _3623_ _3630_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ dacArea_dac_cnt_2\[4\] net13 _3573_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_23_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6280__A1 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5083__A2 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input102_I wb_DAT_MOSI[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6032__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _0301_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ _2548_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3928_ _3461_ _3453_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6647_ _2405_ _2406_ _2411_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3859_ _3399_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6578_ _2412_ _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A2 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _1253_ _1255_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout220 net221 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4337__A1 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5837__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _0744_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5880_ _1631_ _1642_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _0681_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6565__A2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7550_ _0070_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4576__A1 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _0615_ _0461_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6501_ _2298_ _2332_ _2337_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ net74 net73 net76 net75 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7481_ _0001_ net211 dacArea_dac_cnt_3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4693_ _0547_ _3324_ _0471_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6432_ _2265_ _2266_ _2267_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _2194_ _2195_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_143_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5314_ _1141_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6294_ _2013_ _2014_ _2011_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5245_ _0995_ _0555_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ _1020_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_25_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ dacArea_dac_cnt_4\[0\] net26 _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_25_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4058_ _3559_ _3561_ _3562_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6005__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3943__I _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5819__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_240 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_251 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__6492__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_262 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7540__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _0423_ _0879_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _2810_ _2811_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4797__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _1234_ _3396_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_81_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__B _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5863_ _1595_ _1596_ _1594_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6538__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7602_ _0122_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4549__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _0315_ _0462_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5794_ _1636_ _3332_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7533_ _0053_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0598_ _0558_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7464_ _0138_ net203 dacArea_dac_cnt_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4676_ _0474_ _0530_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6415_ dspArea_regP\[24\] _2252_ _1619_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7395_ _0379_ _3216_ _3217_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_1_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6346_ _0327_ _1346_ _2083_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7266__A3 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6277_ _1367_ dspArea_regA\[23\] _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput107 wb_DAT_MOSI[17] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput118 wb_DAT_MOSI[4] net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5228_ _0934_ _1075_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input30_I la_data_in[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__I _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5159_ _0941_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7563__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6701__A2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__A3 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6465__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6768__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A1 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__I _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ _3291_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _0328_ net100 _0316_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7055__I _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6200_ _1821_ _1822_ _1826_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_7180_ _2994_ _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4392_ _0267_ net99 _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1970_ _0956_ _1870_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ dspArea_regP\[21\] _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ _0692_ _0703_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _3481_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1754_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6895_ _0928_ _3449_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5777_ _0882_ _1620_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7516_ _0036_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4728_ _0529_ _0532_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input78_I wb_ADR[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7447_ dspArea_regP\[46\] _0370_ _3255_ _3260_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7378_ _3167_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _2087_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5422__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3984__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6922__A2 _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4499__I _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7459__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ dspArea_regP\[29\] _3420_ net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5964__A3 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _0346_ _3330_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6680_ _2306_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3892_ dspArea_regP\[17\] _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7166__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5177__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _1472_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5793__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6913__A2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4924__A1 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7301_ _3123_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4513_ _0267_ _3301_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ _1316_ _1318_ _1337_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7232_ _3050_ _3058_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4444_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6141__A3 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7163_ _2919_ _2935_ _2990_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4375_ _3469_ _0247_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6429__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _1871_ _1874_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7094_ _2774_ _2776_ _2850_ _2771_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_59_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _0614_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5101__A1 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__C _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A2 _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7157__A2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _2708_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _0465_ _1478_ _1474_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_10_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output184_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6668__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6748__B _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7601__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4143__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5891__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6840__A1 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7396__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6199__A3 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3957__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4906__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4160_ dacArea_dac_cnt_4\[6\] net32 _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_68_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4091_ dacArea_dac_cnt_3\[0\] net17 _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6831__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5634__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__I _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6801_ _2556_ _2564_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_24_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5398__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4993_ _0837_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__A3 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3944_ _3475_ _3453_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6732_ _2553_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6663_ _2483_ _2497_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_143_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3875_ _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6412__I _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6898__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5614_ _0308_ _3361_ _1354_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ _2335_ _2336_ _2332_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ _1387_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4373__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5570__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _0340_ _0920_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7215_ _2249_ _2929_ _3042_ _2928_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__4125__A2 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4427_ _0288_ _0299_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3771__I _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ _2973_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4358_ _0242_ _0238_ _0243_ _0241_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_28_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7077_ _2902_ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4289_ _3294_ _0191_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6822__A1 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6028_ _1022_ _3389_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_73_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4364__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5313__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5616__A2 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3856__I _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5330_ _0897_ _1175_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5261_ _0330_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5304__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7063__I _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7000_ _1190_ _3443_ _2661_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4212_ _3681_ _3683_ _3684_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5192_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ dacArea_dac_cnt_4\[3\] net29 _3629_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6804__A1 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ dacArea_dac_cnt_2\[4\] net13 _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6032__A2 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__A1 dacArea_dac_cnt_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4976_ _0809_ _0813_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6715_ _2463_ _2476_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3927_ _3460_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6646_ _2386_ _2480_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3858_ _3398_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5543__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _2405_ _2406_ _2411_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3789_ _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5528_ _1365_ _1371_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA_input60_I la_data_in[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _1013_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout221 net222 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7048__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output147_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ dspArea_regP\[32\] _2857_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_75_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6023__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5782__A1 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5534__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__A3 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4300__I _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5837__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _0671_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4191__B _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ net79 net78 net81 net80 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_6500_ _2335_ _2336_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7480_ _0000_ net211 dacArea_dac_cnt_3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3784__C2 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4692_ _0283_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _2265_ _2266_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__5525__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6362_ _2196_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5313_ _1157_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6293_ _2013_ _2014_ _2011_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5244_ _1090_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _1021_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _3522_ _3616_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__A1 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4057_ _3557_ _3560_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7202__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7396__C _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4567__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4959_ _0759_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _2301_ _2311_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_4_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5819__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_230 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_241 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_252 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_263 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7492__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__A1 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5886__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7432__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4246__A1 _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _1755_ dspArea_regA\[23\] _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_65_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _0307_ _3391_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4797__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__A1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _1595_ _1596_ _1594_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_34_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7601_ _0121_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _0664_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5746__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _0352_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _0052_ clknet_3_4__leaf_wb_clk_i dspArea_regA\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4744_ _0550_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7463_ _0137_ net201 dacArea_dac_cnt_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4675_ _0481_ _0483_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6414_ _2240_ _2251_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7394_ _3200_ _3202_ _3215_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6345_ _1759_ _3407_ _1965_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6276_ _1149_ _3465_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput108 wb_DAT_MOSI[18] net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5227_ _0971_ _0972_ _0970_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput119 wb_DAT_MOSI[5] net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ _0946_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input23_I la_data_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109_ _3601_ _3599_ _3602_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7423__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A1 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _0465_ _0470_ _0773_ _0834_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_84_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4788__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6162__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6465__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7414__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4779__A2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__I _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4460_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4391_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6130_ _1018_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _0697_ dspArea_regA\[21\] _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5012_ _0845_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_79_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _0309_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5914_ _1755_ _3383_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_81_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _2722_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_62_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _1684_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5195__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5776_ dspArea_regP\[18\] _1618_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7515_ _0035_ net217 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4727_ _0529_ _0532_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3774__I _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7446_ dspArea_regP\[46\] _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6144__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ dspArea_regB\[3\] _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 wb_ADR[31] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7377_ _3189_ _3192_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4589_ _0445_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6328_ _2153_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _0607_ _1884_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3949__I _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7530__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5949__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__I _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__A2 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ dspArea_regP\[28\] _3486_ net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _3411_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_43_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _1473_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_31_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6374__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5177__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4924__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7300_ _3124_ _3125_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ dspArea_regP\[0\] _0267_ _3294_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5492_ _1316_ _1318_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7231_ _3047_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4443_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7162_ _2919_ _2935_ _2990_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_4374_ net113 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6429__A2 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ _1871_ _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _2921_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6044_ _0678_ _1884_ _1786_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7553__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input125_I wb_WE vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3769__I _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _2616_ _2698_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ _2706_ _2707_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_23_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5828_ _1669_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_10_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input90_I wb_ADR[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3718__A3 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ _1494_ _1497_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6117__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6668__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7429_ _3365_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4679__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5891__A3 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7576__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ dacArea_dac_cnt_3\[0\] net17 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6800_ _2630_ _2631_ _2632_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_84_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4992_ _0838_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _2556_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3943_ _3474_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4070__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _2487_ _2492_ _2496_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3874_ dspArea_regA\[16\] _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5613_ _0829_ _3377_ _1236_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _2399_ _2425_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5544_ _1202_ _1388_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5570__A2 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5475_ _0346_ _0670_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7214_ _3041_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4426_ _0298_ net119 _0293_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7145_ _1847_ _3444_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4357_ _3427_ _0235_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7075__A2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7076_ _2904_ _2905_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4288_ _0188_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5086__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4883__I dspArea_regB\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _0815_ _0958_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6586__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _2676_ _2679_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_70_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7599__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5313__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A1 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5838__B _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5001__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6501__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ _0347_ _0461_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _3680_ _3682_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5191_ _0283_ _0278_ _1039_ _3359_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_69_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4142_ dacArea_dac_cnt_4\[2\] net28 _3628_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _3570_ _3574_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6804__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4815__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4208__I _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4043__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _2466_ _2475_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3926_ _3459_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _2391_ _2394_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3857_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6576_ _2405_ _2406_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3788_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _1250_ _1252_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3782__I _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _0342_ _3324_ _1111_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA_input53_I la_data_in[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout200 net201 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4409_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout211 net215 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _0554_ _3366_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xfanout222 net223 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7128_ _2934_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _2803_ _2816_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5502__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6731__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A3 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7039__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5470__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4760_ dspArea_regB\[7\] _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3784__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3711_ net83 net82 net85 net84 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__3784__B2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _0503_ _0510_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1847_ _3378_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6399__B _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _2197_ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ _1056_ _1158_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6292_ _2092_ _2127_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _1006_ _1031_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5174_ _1022_ dspArea_regA\[5\] _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ net196 net25 _3615_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _3557_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6862__B _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7202__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A3 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3777__I _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5764__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4958_ _0739_ _0750_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _3444_ _3418_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4889_ _0680_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6628_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6713__A1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5516__A2 dspArea_regA\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ _2386_ _2391_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__4401__I _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A2 _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_231 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_242 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_59_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_253 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_264 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7441__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6180__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5930_ _0460_ _3408_ _1687_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5861_ _1668_ _1700_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7600_ _0120_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4812_ _0610_ _0620_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5792_ _1634_ _3332_ _1547_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _0051_ clknet_3_6__leaf_wb_clk_i dspArea_regA\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4743_ _0544_ _0595_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7462_ _0136_ net203 dacArea_dac_cnt_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4674_ _0481_ _0483_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6413_ _2246_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7393_ _3200_ _3202_ _3215_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6171__A2 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _2178_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7120__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6275_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput109 wb_DAT_MOSI[19] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5226_ _0971_ _0972_ _0970_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5682__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5157_ _1004_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4108_ dacArea_dac_cnt_3\[3\] net20 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5088_ _0846_ _0848_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5434__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I la_data_in[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _3543_ _3547_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A1 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3970__I _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7178__A1 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6521__I _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7350__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6153__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout203_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _3283_ _3275_ _3279_ _0186_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _0694_ _3448_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I la_data_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5011_ _0857_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6962_ dspArea_regP\[30\] _2713_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5600__I dspArea_regB\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5967__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5913_ _1116_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7169__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6893_ _2723_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5844_ _1685_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5775_ _0395_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7514_ _0034_ net221 dacArea_dac_cnt_7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4726_ _0560_ _0577_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__7482__CLK net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7445_ _0154_ _3259_ _3261_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ _0290_ _0466_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput80 wb_ADR[22] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7376_ dspArea_regP\[39\] _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput91 wb_ADR[3] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4588_ _0398_ _0418_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6327_ _2156_ _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3790__I _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6258_ _0460_ _3434_ _1996_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5209_ dspArea_regA\[13\] _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _1923_ _1926_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5407__A1 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6080__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5666__B _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__I _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6135__A2 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7399__A1 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3890_ _3427_ _3418_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6374__A2 dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5177__A3 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3875__I _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5560_ _1297_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4511_ _0364_ _0372_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7323__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6126__A2 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5491_ _1320_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7230_ _3055_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4442_ dspArea_regB\[8\] _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5885__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7161_ _2938_ _2989_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4373_ _0253_ _0250_ _0254_ _0252_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6200__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _1874_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6429__A3 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7092_ _2616_ _2698_ _2771_ _2850_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1478_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6062__A1 dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input118_I wb_DAT_MOSI[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _2774_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _2706_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ _0307_ _0956_ _1570_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ _1537_ _1598_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_6_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input83_I wb_ADR[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _0282_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5689_ _1197_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7428_ _0426_ _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7359_ _3178_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5800__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6356__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A3 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4520__S _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _0840_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _2562_ _2563_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3942_ _3473_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3802__C2 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _2494_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3873_ _3412_ net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4358__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5612_ _1455_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6592_ _2426_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5543_ _1265_ _1268_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _1228_ _1319_ _1240_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7213_ _2917_ _2918_ _2990_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4425_ _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7520__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7144_ _2971_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4356_ net107 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _2823_ _2839_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4287_ _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5086__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1019_ _3376_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6586__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6928_ _2676_ _2679_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _2681_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4404__I _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5849__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4521__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6274__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6026__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6577__A2 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A2 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7543__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _3680_ _3682_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A1 dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ _3625_ _3627_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__A1 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4072_ dacArea_dac_cnt_2\[4\] net13 _3573_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4815__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A1 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4974_ _0823_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ _2453_ _2454_ _2547_ _2354_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3925_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6644_ _2391_ _2478_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _2407_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3787_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4751__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ dspArea_regP\[15\] _1251_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _1302_ _1220_ _1223_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4503__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout201 net209 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5388_ _1234_ _0949_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout212 net214 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout223 net65 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input46_I la_data_in[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7127_ _2951_ _2955_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4339_ _0226_ _0227_ _0228_ _0229_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_59_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _2886_ _2887_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6009_ _1844_ _1846_ _1848_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__I _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7566__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4990__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6731__A2 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6247__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6970__A2 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _3265_ net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _0488_ _0491_ _0538_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4733__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _1352_ _3438_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _1062_ _1064_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _2128_ _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5289__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ _1010_ _1030_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5173_ _0312_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6238__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ _3613_ _3611_ _3614_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6789__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 la_data_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4055_ dacArea_dac_cnt_2\[1\] net9 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_72_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5461__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7589__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input100_I wb_DAT_MOSI[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _3443_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4972__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ _0666_ _0734_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__I _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3839_ _3280_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6627_ _2370_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6713__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _2392_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _1350_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6489_ _2318_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_232 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_243 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_254 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_59_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XDSP48_265 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__A3 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5452__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3968__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4963__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6519__I dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5443__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3878__I _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _1701_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _0663_ _0619_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _0348_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4742_ _0590_ _0592_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_7530_ _0050_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7461_ _0135_ net200 dacArea_dac_cnt_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4673_ _0520_ _0524_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4502__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7392_ _3213_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6343_ _2179_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6274_ _2107_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7120__A2 _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _1032_ _1070_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_69_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5682__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5156_ _0917_ _0931_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ dacArea_dac_cnt_3\[3\] net20 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_29_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5087_ _0935_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ dacArea_dac_cnt_1\[5\] net5 _3546_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4493__I0 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5985__A3 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7187__A2 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ dspArea_regP\[21\] _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7659_ net197 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7604__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7111__A2 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 wb_DAT_MISO[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3987__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A3 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7350__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A1 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _0858_ _0859_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__A1 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6961_ _2763_ _2766_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _0736_ _0955_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_46_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7169__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _1110_ _3439_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7413__I0 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ dspArea_regB\[2\] dspArea_regA\[17\] _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5774_ _1610_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6392__A3 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7513_ _0033_ net220 dacArea_dac_cnt_7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4725_ _0520_ _0578_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7444_ _0425_ _3247_ _3252_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_4656_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7341__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput70 wb_ADR[13] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput81 wb_ADR[23] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5352__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _0413_ _0417_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7375_ _0495_ _3197_ _3198_ _3521_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput92 wb_ADR[4] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6326_ _2162_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_1_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _0285_ _3450_ _1898_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6852__A1 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _0570_ _3384_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6188_ _1923_ _1926_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5139_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__I dspArea_regB\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4918__A1 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5591__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__I _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4146__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ dspArea_regP\[0\] _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_8_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _1326_ _1331_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7323__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5334__A1 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _0163_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3891__I _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7160_ _2985_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4372_ _3461_ _0247_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1938_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _2239_ _2348_ _2441_ _2542_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _0675_ _3433_ _1686_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6062__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _2700_ _2701_ _2615_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__4073__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ _0760_ _3473_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ _0302_ _3391_ _1465_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4376__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _1457_ _1599_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4708_ _0562_ _3315_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7314__A2 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _1530_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input76_I wb_ADR[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ _3225_ _3244_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_68_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5325__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ dspArea_regP\[5\] _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7358_ _3179_ _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_11_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _3498_ _2044_ _2147_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_7289_ _0360_ _3461_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__I0 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5521__I dspArea_regB\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__I0 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5800__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4119__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A2 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7241__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6044__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4990_ _0296_ _3335_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _3472_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3802__B2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3872_ dspArea_regP\[47\] _3382_ _3310_ _3410_ _3411_ dspArea_regP\[15\] _3412_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6660_ _1450_ _3415_ _2390_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _1430_ _1432_ _1454_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6591_ _2312_ _2331_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5542_ _1265_ _1268_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5307__A1 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _1230_ _1231_ _1238_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7212_ _2919_ _3039_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4424_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4355_ _0237_ _0238_ _0239_ _0241_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7143_ _1416_ _3443_ _2867_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_59_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6807__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7074_ _2903_ _2822_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _0188_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6025_ _1862_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4294__A1 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4046__A1 dacArea_dac_cnt_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _2746_ _2758_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4597__A2 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3796__I _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _2684_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_13_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _0339_ _3343_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5546__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _2239_ _2348_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7495__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6274__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A1 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4512__A2 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4140_ dacArea_dac_cnt_4\[2\] net28 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _3571_ _3568_ _3572_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_23_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4276__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A2 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__A1 _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4973_ _0335_ _3292_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6712_ _0423_ _2545_ _2546_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3924_ _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6643_ _2394_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3855_ _3395_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6574_ _2408_ _2409_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3786_ dspArea_regA\[6\] _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__A3 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5525_ _1366_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4751__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5456_ _1139_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4407_ dspArea_regB\[3\] _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5700__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout202 net209 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout213 net214 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2952_ _2954_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4338_ _0193_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input39_I la_data_in[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4269_ _0173_ _0174_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7057_ _2835_ _2836_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6008_ _1844_ _1846_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_68_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4019__A1 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A3 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__I dspArea_regB\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7444__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__A2 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5758__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4325__I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7510__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__I _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5930__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _1062_ _1064_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6290_ _1991_ _2010_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5241_ _0824_ _0997_ _1001_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5172_ _0319_ _0920_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ dacArea_dac_cnt_3\[6\] net24 _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6238__A2 dspArea_regA\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4054_ _3558_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 la_data_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _0744_ _0751_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3907_ _3442_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _0602_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6626_ _1297_ _3379_ _2371_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3838_ _3381_ net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6557_ _0326_ _3406_ _2289_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5921__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _3280_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5508_ _1351_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6488_ _2321_ _2324_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _1184_ _1281_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_233 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_244 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_255 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_19_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_266 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_output145_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7109_ _2936_ _2937_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5988__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7533__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4660__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6401__A2 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7417__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4810_ _0613_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5790_ _1632_ _3347_ _1439_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4741_ _0590_ _0592_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3894__I dspArea_regA\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _0134_ net200 dacArea_dac_cnt_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4672_ _0525_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _1509_ _1510_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5903__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ _3210_ _3212_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6951__I0 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6342_ _0313_ _3413_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6273_ _2109_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5224_ _1071_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5131__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _0923_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_5_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6873__C _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4106_ _3596_ _3600_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5086_ _0838_ _0842_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ _3544_ _3545_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_65_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__I1 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7187__A3 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6395__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _0882_ _1829_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4939_ _0710_ _0711_ _0709_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7658_ net198 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6609_ _2150_ _2234_ _2347_ _2255_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7589_ _0109_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput180 net180 wb_DAT_MISO[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput191 net191 wb_DAT_MISO[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__I _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7598__D _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4603__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A2 dspArea_regA\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7579__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3889__I _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__A2 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6960_ _2789_ _2790_ _2762_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_35_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ _0326_ _3367_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_35_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6891_ _0996_ _1992_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A1 dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5842_ dspArea_regB\[3\] _1368_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5773_ _1292_ _1611_ _1613_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_33_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7512_ _0032_ net218 dacArea_dac_cnt_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4724_ _0524_ _0528_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6129__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7443_ dspArea_regP\[45\] dspArea_regP\[44\] _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4655_ _0503_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 la_data_in[63] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7374_ dspArea_regP\[38\] _0426_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput71 wb_ADR[14] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5352__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput82 wb_ADR[24] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4586_ _0410_ _0439_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xinput93 wb_ADR[5] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6325_ _1533_ _3363_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6256_ _2093_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5207_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _1936_ _2021_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_5138_ _0367_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_40_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input21_I la_data_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3799__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _0815_ _3312_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__I _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5591__A2 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4606__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6359__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5582__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4440_ _0288_ _0310_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5334__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ net112 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5164__I _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6110_ _1941_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ _2917_ _2919_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1880_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4508__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _2630_ _2631_ _2697_ _2632_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_23_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6874_ _0828_ _3480_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _1666_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4243__I _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5756_ _1491_ _1492_ _1490_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6770__A1 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4707_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ _1526_ _1528_ _1529_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7426_ _3238_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4638_ _0425_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input69_I wb_ADR[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7357_ _3180_ _3151_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4569_ _0279_ _3305_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5074__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6308_ _2045_ _2145_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7288_ _3112_ _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5089__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _2076_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5802__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4687__I1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4418__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4439__I1 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6761__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4328__I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6044__A3 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ dspArea_regA\[23\] _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3871_ _3295_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5004__A1 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _1430_ _1432_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__6752__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _2326_ _2330_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5555__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5541_ _1314_ _1383_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _1211_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7211_ _2938_ _2989_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4423_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7142_ _1414_ _3459_ _2806_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4354_ _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6807__A2 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7073_ _2819_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4285_ _0187_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4818__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _1863_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_39_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4294__A2 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input123_I wb_DAT_MOSI[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _2750_ _2757_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_70_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5794__A2 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _2688_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _1435_ _0769_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _2620_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5739_ _1150_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_13_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7409_ _3199_ _3148_ _2795_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_11_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6628__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4809__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5482__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6982__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__I dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A3 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4070_ dacArea_dac_cnt_2\[3\] net11 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5473__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3897__I _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _0819_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_63_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__A1 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6711_ _2542_ _2544_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3923_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6642_ _2463_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3854_ dspArea_regA\[14\] _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6573_ _1134_ dspArea_regA\[21\] _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3785_ _3334_ net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4200__A2 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ dspArea_regP\[16\] _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5455_ _1129_ _1140_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4406_ _0262_ _0281_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5386_ dspArea_regB\[6\] _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5700__A2 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout203 net208 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_5_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7125_ _2868_ _2953_ _2952_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4337_ _3387_ _0224_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7056_ _2885_ _2834_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4268_ dacArea_dac_cnt_7\[4\] net57 _0171_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__A2 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6007_ _1847_ _3347_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4199_ _3666_ _3674_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7205__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5767__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6909_ _2652_ _2674_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7462__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5262__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7444__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4194__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout219_I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A2 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7132__A1 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7652__I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _1079_ _1081_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_5_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5171_ _1019_ _0670_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ dacArea_dac_cnt_3\[6\] net24 _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4053_ _3487_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput3 la_data_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6946__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _0802_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6410__A3 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3906_ _3441_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4886_ _0737_ _3299_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7485__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _2458_ _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3837_ dspArea_regP\[43\] _3351_ _3373_ _3379_ _3380_ dspArea_regP\[11\] _3381_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__7371__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _0321_ _1582_ _2180_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_69_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3768_ _3319_ net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5921__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ _1352_ _0955_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6487_ _2211_ _2213_ _2323_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ _1082_ _1176_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input51_I la_data_in[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ _1212_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_234 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_245 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_256 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_7108_ _2907_ _2911_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XDSP48_267 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_47_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7039_ _0737_ _2210_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6165__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5912__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4537__S _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4100__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__I _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _0497_ _0594_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ dspArea_regP\[6\] _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7353__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _2247_ _1824_ _2039_ _2241_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7390_ _3210_ _3212_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6951__I1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6341_ _0815_ _3404_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _0468_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _0948_ _0969_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5154_ _0930_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4105_ dacArea_dac_cnt_3\[3\] net20 _3599_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_29_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ _0303_ _3339_ _0763_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4036_ dacArea_dac_cnt_1\[4\] net4 _3541_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_53_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6919__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ dspArea_regP\[20\] _1828_ _1619_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ _0710_ _0711_ _0709_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input99_I wb_DAT_MOSI[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7657_ net199 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7344__A1 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _0717_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5077__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ _2256_ _2442_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7588_ _0108_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _2362_ _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput170 net170 wb_DAT_MISO[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput181 net181 wb_DAT_MISO[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7500__CLK net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6083__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6138__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6689__A3 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5649__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A2 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6861__A3 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5821__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ _1748_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _0347_ _3424_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _0622_ _3405_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6377__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5772_ _1401_ _1614_ _1615_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_21_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7511_ _0031_ net220 dacArea_dac_cnt_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4723_ _0524_ _0528_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7326__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7442_ dspArea_regP\[45\] _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4654_ _0506_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
Xinput50 la_data_in[54] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7373_ _3193_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xinput61 la_data_in[6] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput72 wb_ADR[15] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4585_ _0440_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput83 wb_ADR[25] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput94 wb_ADR[6] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7523__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6324_ _2160_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_66_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _0608_ _3409_ _1986_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6301__A2 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _1051_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6186_ _2024_ _2025_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_57_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5137_ net125 _3276_ _0365_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6065__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _0747_ _0466_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input14_I la_data_in[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4019_ _3489_ _3530_ _3531_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_53_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4551__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6056__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4606__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6359__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7546__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6531__A2 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout201_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _0249_ _0250_ _0251_ _0252_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7660__I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _0308_ _1346_ _1777_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I la_data_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A2 dspArea_regA\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6047__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6598__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _2633_ _2772_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_35_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6873_ _0988_ _2704_ _2705_ _2354_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5824_ _1646_ _1648_ _1665_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ _1491_ _1492_ _1490_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_31_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _0289_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5686_ _1526_ _1528_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_8_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ _0452_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7425_ _3240_ _3237_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7356_ _3150_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4568_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6307_ _2140_ _2144_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7287_ _3109_ _3110_ _3111_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4499_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5089__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _1109_ dspArea_regA\[12\] _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _2006_ _2007_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6589__A2 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4434__I dspArea_regB\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7569__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6210__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6761__A2 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__A1 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6277__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4609__I _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5004__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7655__I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _1224_ _1384_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5471_ _1216_ _1219_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7210_ _2938_ _2989_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4515__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ dspArea_regB\[5\] _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7141_ _2967_ _2968_ _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4353_ net126 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6268__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7072_ _2884_ _2901_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4284_ _3278_ _3285_ _0186_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4818__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6023_ _0331_ _1038_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4519__I _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input116_I wb_DAT_MOSI[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ _2755_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _1198_ _3401_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ _1564_ _1649_ _1573_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_13_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3999_ _3488_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6787_ _2457_ _2541_ _2437_ _2440_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_50_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5738_ _3422_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I wb_ADR[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _0989_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4506__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _0362_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7339_ _3163_ _3117_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_output168_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6259__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4809__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6982__A2 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4993__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6734__A2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3720__A2 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout199_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6670__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _0820_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6973__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6710_ _2542_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3922_ dspArea_regA\[21\] _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4984__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ _3394_ net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6641_ _2466_ _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6725__A2 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ dspArea_regP\[37\] _3320_ _3311_ _3333_ _3318_ dspArea_regP\[5\] _3334_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6572_ _1233_ _2108_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5523_ _1367_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6489__A1 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5454_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _0280_ net116 _0269_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5385_ _0307_ _3354_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout204 net208 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4336_ _0215_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7124_ _2875_ _2876_ _2873_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout215 net222 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _2833_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4267_ dacArea_dac_cnt_7\[4\] net57 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6006_ _1418_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6661__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4198_ dacArea_dac_cnt_5\[6\] net41 _3673_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_27_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__A1 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _2738_ _2739_ _2651_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _2668_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4718__A1 dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6891__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5170_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4121_ _3596_ _3612_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _3492_ _3556_ _3557_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_68_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 la_data_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7199__A2 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _0803_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6410__A4 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3905_ _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6624_ _2362_ _2374_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3836_ _3296_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3767_ dspArea_regP\[35\] _3281_ _3311_ _3317_ _3318_ dspArea_regP\[3\] _3319_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6555_ _2387_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5921__A3 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5506_ _0295_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6486_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5437_ _1174_ _1274_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6882__A1 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _1213_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XDSP48_224 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_235 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_input44_I la_data_in[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_246 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_7107_ _2902_ _2906_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XDSP48_257 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_4319_ net122 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5299_ _1142_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_87_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7038_ _2864_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_68_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4707__I _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4442__I dspArea_regB\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A3 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5373__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__I0 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5987__I0 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _0265_ _3337_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7353__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _0747_ _3397_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_31_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6271_ dspArea_regA\[21\] _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _0965_ _0968_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _0998_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4104_ dacArea_dac_cnt_3\[2\] net19 _3598_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6616__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5084_ _0909_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ dacArea_dac_cnt_1\[4\] net4 _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7452__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__A2 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7041__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1818_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_12_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4937_ _0752_ _0785_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_7656_ net192 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _0719_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7344__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _2259_ _2438_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3819_ _3364_ net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7587_ _0107_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4799_ _0586_ _0589_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ _2365_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _1134_ _3447_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6855__A1 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput160 net160 wb_DAT_MISO[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput171 net171 wb_DAT_MISO[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output150_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput182 net182 wb_DAT_MISO[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4469__I0 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__I _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5830__A2 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5594__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__I dspArea_regB\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5346__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7099__A1 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4347__I _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7658__I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _1671_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_62_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5771_ _1404_ _1607_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7510_ _0030_ net220 dacArea_dac_cnt_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _0569_ _0574_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_33_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__A2 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__A3 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ dspArea_regP\[44\] _0425_ _3247_ _3252_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__5337__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _0457_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput40 la_data_in[45] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4810__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput51 la_data_in[55] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7372_ _3167_ _3195_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput62 la_data_in[7] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4584_ _0406_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput73 wb_ADR[16] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput84 wb_ADR[26] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 wb_ADR[7] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6323_ _2157_ _2158_ _2159_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _0829_ _3426_ _1889_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_66_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5205_ _1052_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6185_ _1855_ _1922_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5136_ _3271_ _3277_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _0914_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ _3528_ _3529_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__A2 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4379__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5969_ _1644_ _1708_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5879__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6828__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7498__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4303__A2 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4067__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7005__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A3 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7308__A2 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6531__A3 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4542__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6047__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A1 _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6941_ _2636_ _2768_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_19_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ dspArea_regP\[29\] _0380_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_62_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _1646_ _1648_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_37_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5754_ _1561_ _1594_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _0509_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5685_ _1418_ _3325_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _3233_ _3239_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4636_ _0453_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7355_ _0356_ _3149_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4533__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _3287_ _0368_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6306_ _2140_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7286_ _3109_ _3110_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4498_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5089__A3 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _1437_ _3374_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4297__A1 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _1904_ _1906_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _0965_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4049__A1 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _1770_ _1781_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5797__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5320__B _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__I _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6210__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4221__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4450__I _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6277__A2 dspArea_regA\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7226__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7513__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4561__S _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6201__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4212__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5470_ _1216_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4421_ _0288_ _0294_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4515__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7671__I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7140_ _2859_ _2878_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4352_ _3417_ _0235_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6268__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7071_ _2888_ _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4283_ net98 net125 net159 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6022_ _0340_ _3358_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6951__S _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _1424_ _3409_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6440__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input109_I wb_DAT_MOSI[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6855_ _2686_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5806_ _1565_ _1566_ _1571_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4203__A1 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _2457_ _2541_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3998_ _3499_ _3514_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5737_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5668_ _1504_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input74_I wb_ADR[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4506__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _0263_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5599_ _1443_ _1045_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7338_ _3106_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6259__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7269_ _3037_ _3086_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7536__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4445__I _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__A2 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5942__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__A1 dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__C _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _0748_ _0552_ _0746_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _3454_ _3455_ net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4984__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7666__I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _2473_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3852_ dspArea_regP\[45\] _3382_ _3373_ _3393_ _3380_ dspArea_regP\[13\] _3394_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6571_ _0614_ _3440_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3783_ _3332_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5522_ dspArea_regA\[16\] _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5453_ _1195_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5384_ _0460_ _3369_ _1146_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7438__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7123_ _2875_ _2876_ _2873_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout205 net207 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4335_ net102 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7559__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout216 net218 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7054_ _2880_ _2883_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6110__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4266_ _0164_ _0172_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_45_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6005_ _1845_ _3347_ _1751_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_86_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6661__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ dacArea_dac_cnt_5\[5\] net40 _3672_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_28_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6413__A2 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _2638_ _2647_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _2596_ _2669_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_51_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5924__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6769_ _2585_ _2589_ _2602_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7429__A1 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6340__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4120_ dacArea_dac_cnt_3\[6\] net24 _3611_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4051_ dacArea_dac_cnt_2\[0\] net8 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 la_data_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _0729_ _0795_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3904_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7672_ net192 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6159__A1 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4884_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6623_ _2365_ _2373_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3835_ _3378_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5906__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6554_ _2388_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3766_ _3296_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _0839_ _1039_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ dspArea_regP\[24\] _0265_ _2319_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _1184_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6331__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ _0312_ dspArea_regA\[7\] _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_225 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4893__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_236 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_7106_ _2920_ _2931_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XDSP48_247 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_4318_ _0211_ _0204_ _0213_ _0206_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XDSP48_258 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5298_ _1143_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input37_I la_data_in[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ _2865_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6634__A2 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4249_ _0156_ _0157_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__I1 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6873__A2 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7050__A2 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5987__I1 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5061__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7165__B _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6313__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _0515_ _2108_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _1050_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _0999_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _3594_ _3597_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6616__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5419__A3 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _0913_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4627__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4034_ _3515_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__A2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5985_ _1821_ _1822_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4936_ _0786_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_36_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ net193 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _0654_ _0652_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6606_ _2259_ _2438_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3818_ dspArea_regP\[41\] _3351_ _3342_ _3363_ _3349_ dspArea_regP\[9\] _3364_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7586_ _0106_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6552__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _0648_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_20_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _2371_ _2372_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3749_ dspArea_regP\[33\] _3281_ _3289_ _3302_ _3297_ dspArea_regP\[1\] _3303_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5107__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _1233_ _3438_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5419_ _1163_ _1164_ _1162_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5658__A3 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput150 net150 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput161 net161 wb_DAT_MISO[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6399_ _2136_ _2137_ _2135_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput172 net172 wb_DAT_MISO[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput183 net183 wb_DAT_MISO[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__B _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output143_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4618__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__I1 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__I _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__A1 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5594__A2 dspArea_regA\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6543__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7099__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5821__A3 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4363__I _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _1404_ _1607_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4721_ _0525_ _0527_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7440_ _3492_ _3257_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _0507_ dspArea_regA\[1\] _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput30 la_data_in[36] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7371_ _3133_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput41 la_data_in[46] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput52 la_data_in[56] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4583_ _0411_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput63 la_data_in[8] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput74 wb_ADR[17] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6322_ _2157_ _2158_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
Xinput85 wb_ADR[27] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput96 wb_ADR[8] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4739__S _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6253_ _2090_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4848__A1 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5204_ _0277_ _0955_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6184_ _1919_ _2023_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5135_ _0882_ _0984_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5066_ _0915_ _0552_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5273__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _3528_ _3529_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_84_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6773__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5968_ _1704_ _1707_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_40_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4919_ _0470_ _3353_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5899_ _1728_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7569_ _0089_ clknet_3_3__leaf_wb_clk_i dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6828__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6149__B _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5264__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7005__A2 _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__A3 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__A1 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7592__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7669__I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6940_ _2636_ _2768_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _2698_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5189__I dspArea_regA\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ _1650_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5753_ _1595_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5917__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _0550_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _1527_ _3325_ _1440_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_72_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7423_ _0988_ _3242_ _3243_ _3521_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4635_ _0488_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _3176_ _3177_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6305_ _2141_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7285_ _0354_ _3468_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4497_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6236_ _1435_ _1039_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5089__A4 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4297__A2 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _1904_ _1906_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _0850_ _0966_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_57_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1850_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_73_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _0869_ _0872_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5099__I dspArea_regA\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7465__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A2 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__I _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5562__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7226__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5237__A1 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _0292_ net118 _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3723__A1 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _0215_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7070_ _2891_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4282_ net99 _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5476__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _1012_ _3353_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _2753_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_82_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6854_ _0353_ _3409_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_39_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7488__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5805_ _1548_ _1647_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_17_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6785_ _2444_ _2446_ _2617_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3997_ dacArea_dac_cnt_0\[5\] net56 _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4203__A2 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5736_ _1576_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__A1 dspArea_regP\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5667_ _1506_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7406_ _3226_ _3227_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4618_ _0273_ _0433_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6900__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ dspArea_regB\[9\] _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input67_I wb_ADR[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7337_ _3108_ _3116_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4549_ _0286_ _3293_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__I _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7268_ _2918_ _3038_ _3039_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_78_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6219_ _2057_ _1973_ _1976_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7199_ _2961_ _2979_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7258__B _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3953__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3805__I dspArea_regA\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7447__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6407__B1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ dspArea_regP\[20\] _3429_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4984__A3 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ _3392_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7383__A1 dspArea_regP\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _0562_ _3458_ _2317_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3782_ _3331_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3944__A1 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ dspArea_regB\[0\] _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _1297_ _0391_ _1196_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__A1 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5383_ _0675_ _1229_ _1053_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_7122_ _2945_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4334_ _0223_ _0216_ _0225_ _0218_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xfanout206 net207 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout217 net218 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_7053_ _2881_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4265_ dacArea_dac_cnt_7\[4\] net57 _0171_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6110__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4121__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _0348_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4196_ _3671_ _3669_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input121_I wb_DAT_MOSI[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _2638_ _2647_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_39_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _2490_ _2665_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7374__A1 dspArea_regP\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4188__A1 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6768_ _2594_ _2598_ _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5924__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _1342_ _3369_ _1466_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6699_ _2426_ _2427_ _2425_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6168__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5915__A2 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7117__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6340__A2 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ dacArea_dac_cnt_2\[0\] net8 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_49_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5851__A1 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 la_data_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _0730_ _0801_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_64_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3903_ _3438_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7671_ net193 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__A2 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ dspArea_regB\[9\] _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _2359_ _2455_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3834_ _3377_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5906__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6553_ _0312_ dspArea_regA\[18\] _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3765_ _3316_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7526__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ _0551_ _0773_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6484_ _2254_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _1273_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__A2 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _0318_ dspArea_regA\[6\] _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XDSP48_226 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__A2 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XDSP48_237 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7105_ dspArea_regP\[33\] _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4317_ _3348_ _0212_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XDSP48_248 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5297_ _1144_ _0958_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XDSP48_259 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7036_ _0332_ _3457_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4248_ _0156_ _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6634__A3 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 dspArea_regB\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ dacArea_dac_cnt_5\[2\] net37 _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7347__A1 _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__A3 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7549__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout217_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7165__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4572__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6313__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _1065_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ _0909_ _0933_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4102_ dacArea_dac_cnt_3\[2\] net19 _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5082_ _0917_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5824__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _3516_ _3542_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4824__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1287_ _1291_ _1611_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_80_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4935_ _0686_ _0708_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7654_ net194 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4866_ _0718_ _0651_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6605_ _2437_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3817_ _3362_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7585_ _0105_ clknet_3_4__leaf_wb_clk_i dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4797_ _0503_ _0510_ _0585_ _0650_ _0581_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__6552__A2 dspArea_regA\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3748_ _3301_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6536_ _1533_ _3379_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _0306_ _3432_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6304__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput140 net140 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5418_ _1224_ _1261_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xoutput151 net151 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6398_ _2136_ _2137_ _2135_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput162 net162 wb_DAT_MISO[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4866__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput173 net173 wb_DAT_MISO[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput184 net184 wb_DAT_MISO[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5349_ _1194_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4618__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5815__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _2848_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_47_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6791__A2 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6059__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5282__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__I _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4720_ dspArea_regP\[6\] _0526_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4651_ dspArea_regB\[6\] _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 la_data_in[27] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 la_data_in[37] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4545__A1 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7370_ _3139_ _3168_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4582_ _0403_ _0405_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput42 la_data_in[47] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput53 la_data_in[57] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput64 la_data_in[9] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput75 wb_ADR[18] net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6321_ _1636_ _3370_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 wb_ADR[28] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_66_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput97 wb_ADR[9] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6252_ _2070_ _2072_ _2089_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4848__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5203_ _0515_ _3366_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6183_ _1920_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5134_ dspArea_regP\[12\] _0983_ _0726_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ _0341_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4016_ dacArea_dac_cnt_1\[1\] net64 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5273__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6222__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5967_ _1741_ _1805_ _1808_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4918_ _0768_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ _1731_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_16_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input97_I wb_ADR[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _0632_ _0634_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7568_ _0088_ clknet_3_3__leaf_wb_clk_i dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6519_ dspArea_regP\[26\] _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7325__I1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7499_ _0019_ net214 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4839__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7105__I dspArea_regP\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__I _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6516__A2 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3808__I _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__A3 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _2699_ _2626_ _2702_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_35_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5821_ _1655_ _1660_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_22_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4766__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5752_ _1471_ _1489_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4703_ _0553_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_30_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5683_ _1013_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6507__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7422_ dspArea_regP\[41\] _0380_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4634_ _0410_ _0489_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_15_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7353_ _0360_ _3475_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4565_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5191__A1 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6304_ _2038_ _2040_ _2142_ _2141_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7284_ _2893_ _3468_ _3054_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4496_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6235_ _1980_ _2073_ _1989_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6691__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6166_ _1900_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _0854_ _0856_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6097_ _1407_ _3340_ _1851_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6443__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _0873_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I la_data_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6713__B _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6999_ _2828_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_40_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4757__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4509__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6004__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3980__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5721__A3 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4459__I _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5237__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4748__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ net106 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3723__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4369__I _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _3645_ _0184_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_3_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6673__A1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6020_ _1770_ _1860_ _1780_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I la_data_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6425__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _1419_ _3417_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4987__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6853_ _2485_ _2660_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _1553_ _1556_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6784_ _2437_ _2440_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3996_ _3511_ _3512_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5735_ _1577_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3962__A2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _1509_ _1510_ _1396_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7405_ _3203_ _3209_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4617_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6900__A2 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ _0325_ _3344_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7336_ _3156_ _3160_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4911__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _0280_ _3301_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7267_ _2249_ _2929_ _3092_ _2928_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4479_ _0343_ net102 _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _1893_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7198_ _2957_ _3025_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _1981_ _1982_ _1987_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4690__A3 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7582__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3953__A2 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5458__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__I dspArea_regA\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__A4 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ _3391_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7383__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4197__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3781_ _3330_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5520_ _0271_ _3406_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _0358_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _0277_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5382_ _3385_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7121_ _2946_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ _3379_ _0224_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout207 net208 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_5_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6646__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout218 net221 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4264_ _0169_ _0167_ _0170_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7052_ _2798_ _2818_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _1414_ _3362_ _1653_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4195_ dacArea_dac_cnt_5\[5\] net40 _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7455__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__A1 _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6949__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7071__A1 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input114_I wb_DAT_MOSI[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6905_ _2717_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _2595_ _2597_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7374__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5385__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4432__I0 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _2599_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3979_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _1033_ _1229_ _1353_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ _2426_ _2427_ _2425_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7094__B _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5649_ _1457_ _1490_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__3906__I _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7319_ dspArea_regP\[36\] _3102_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4360__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4472__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3816__I _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7478__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout197_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput7 la_data_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _0731_ _0732_ _0794_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4382__I _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3902_ dspArea_regA\[19\] _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7670_ net194 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4882_ _0667_ _0668_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _2434_ _2435_ _2433_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5367__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3833_ _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6552_ _0318_ dspArea_regA\[17\] _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3764_ _3315_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5503_ _1348_ _3377_ _1247_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__3726__I _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _1149_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5434_ _3681_ _1181_ _1280_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5365_ _0926_ _0478_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _2856_ _2933_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XDSP48_227 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_4316_ _0200_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDSP48_238 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XDSP48_249 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5296_ dspArea_regB\[2\] _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7035_ _0996_ _3449_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4247_ dacArea_dac_cnt_7\[1\] net53 _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _3639_ _3657_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4493__S _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6398__A3 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _2648_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__I0 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__A1 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7283__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7035__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5597__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _0913_ _0932_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7274__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4101_ _3515_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ _0923_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4088__A1 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4032_ dacArea_dac_cnt_1\[4\] net4 _3541_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5824__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4934_ _0704_ _0707_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_80_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7653_ net195 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _0603_ _0647_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_32_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4840__I _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _2259_ _2438_ _2439_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3816_ _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7584_ _0104_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4012__A1 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _0583_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ _2369_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3747_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6466_ _0562_ _3450_ _2208_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5417_ _1262_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput130 net130 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput141 net141 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6397_ _2150_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput152 net152 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput163 net163 wb_DAT_MISO[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput174 net174 wb_DAT_MISO[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5348_ _1191_ _1192_ _1193_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input42_I la_data_in[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput185 net185 wb_DAT_MISO[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__I _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6068__A2 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5279_ _1033_ _3354_ _0944_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_29_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _2791_ _2792_ _2847_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5815__A2 dspArea_regA\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4874__I0 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7099__A4 _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__A3 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7516__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6782__A3 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4793__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _0504_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xinput10 la_data_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput21 la_data_in[28] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput32 la_data_in[38] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _0431_ _0436_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
Xinput43 la_data_in[48] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput54 la_data_in[58] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6320_ _1527_ _3370_ _2078_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
Xinput65 user_clock2 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput76 wb_ADR[19] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput87 wb_ADR[29] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput98 wb_CYC net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6251_ _2070_ _2072_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_143_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5202_ _0624_ _0773_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6182_ _1767_ _1804_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _0897_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5064_ _0333_ _0462_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _3492_ _3527_ _3528_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5273__A3 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _1668_ _1806_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4917_ _3336_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5981__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _1737_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4848_ dspArea_regP\[8\] _0633_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7567_ _0087_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5733__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _0264_ _3352_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ _2254_ _0424_ _2353_ _2354_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _0018_ net217 dacArea_dac_cnt_5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _0927_ _3406_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3914__I _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__S _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7539__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7410__A1 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6764__A3 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5724__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3824__I _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7229__A1 _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5820_ _1661_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5751_ _1485_ _1488_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6091__B _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4702_ _0508_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5682_ _1413_ _3338_ _1324_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_7421_ _3239_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4633_ _0440_ _0442_ _0439_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5715__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7352_ _0356_ _3483_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4564_ _3288_ _0368_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5191__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6303_ _2027_ _2030_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7283_ _0335_ _3481_ _3052_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4495_ dspArea_regB\[15\] _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6234_ _1981_ _1982_ _1987_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6165_ _1998_ _2002_ _2004_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0854_ _0856_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6096_ _1933_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4565__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5047_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ _2720_ _2735_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6713__C _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _1788_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4757__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5706__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6131__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4693__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6434__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__I _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5239__C _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4920__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7026__I _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ net192 net60 _0183_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_4_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6673__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4385__I dspArea_regB\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6921_ _2751_ _2752_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_35_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6852_ _2590_ _2593_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5803_ _1553_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6783_ _2457_ _2541_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5936__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ dacArea_dac_cnt_0\[4\] net45 _3509_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _1144_ _1368_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _0892_ _0895_ _1175_ _1508_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7404_ _3205_ _3208_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4616_ _0463_ _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5596_ _1436_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7335_ _3157_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4547_ _0403_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4911__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7266_ _3037_ _3041_ _3086_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_1_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6113__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _0268_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6217_ _1882_ _1894_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7197_ _2960_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6148_ _1981_ _1982_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _1800_ _1803_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__I _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4902__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6655__A2 dspArea_regA\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A2 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5091__A1 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3780_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5450_ _1293_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5381_ _1226_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7120_ _2947_ _2948_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4332_ _0200_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net209 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7051_ _2793_ _2797_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
Xfanout219 net220 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4263_ dacArea_dac_cnt_7\[3\] net55 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4657__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _1842_ _1763_ _1766_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4194_ _3666_ _3670_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_41_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5082__A1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _2720_ _2735_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input107_I wb_DAT_MOSI[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6835_ _2664_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6582__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _0748_ _3426_ _2491_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5385__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ _3488_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4432__I1 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ _1559_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6697_ _2501_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5137__A2 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6334__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ _1491_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input72_I wb_ADR[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _0358_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _3123_ _3126_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _3059_ _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_46_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output159_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3922__I dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4753__I _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5584__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A1 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3832__I _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput8 la_data_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_64_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6364__B _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _0731_ _0732_ _0794_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_52_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3901_ _3436_ _3437_ net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_17_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ _0731_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6620_ _2434_ _2435_ _2433_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3832_ _3375_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5367__A2 dspArea_regA\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _0926_ _3414_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3763_ _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5502_ _0677_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6482_ dspArea_regA\[24\] _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6316__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _0989_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5364_ _1207_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7103_ dspArea_regP\[32\] _2932_ _2628_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ net121 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XDSP48_228 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _0514_ _3374_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XDSP48_239 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_59_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _0348_ _3441_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4246_ _0154_ _0155_ _0156_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_45_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4177_ dacArea_dac_cnt_5\[2\] net37 _3656_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__7572__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7044__A2 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _2649_ _2576_ _2650_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5358__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__I1 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3917__I _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7536__D _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6749_ _2494_ _2495_ _2492_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4030__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6858__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5294__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6963__I _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7035__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__I _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4483__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__I dspArea_regB\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7595__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _3570_ _3595_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _0925_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5285__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ _3539_ _3537_ _3540_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1717_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_52_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _0767_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_61_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4260__A2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7652_ net196 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4864_ _0662_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6603_ _2343_ _2346_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3815_ _3360_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7583_ _0103_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4795_ _0511_ _0533_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ _2366_ _2367_ _2368_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _0547_ _3466_ _2111_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5416_ _1141_ _1161_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
Xoutput131 net131 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6396_ _2230_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
Xoutput142 net142 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput153 net153 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4568__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput164 net164 wb_DAT_MISO[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5347_ _1191_ _1192_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput175 net175 wb_DAT_MISO[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput186 net186 wb_DAT_MISO[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7265__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5278_ _1103_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4079__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input35_I la_data_in[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7017_ _2791_ _2792_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_4229_ dacArea_dac_cnt_6\[4\] net48 _3695_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4874__I1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5028__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6776__A1 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4251__A2 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7468__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4478__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5267__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__A3 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout222_I net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput11 la_data_in[19] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput22 la_data_in[29] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4580_ _0399_ _0402_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput33 la_data_in[39] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput44 la_data_in[49] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput55 la_data_in[59] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput66 wb_ADR[0] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput77 wb_ADR[1] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput88 wb_ADR[2] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput99 wb_DAT_MOSI[0] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6250_ _2074_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6089__B _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5201_ _1036_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4388__I _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6181_ _1951_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5132_ _0980_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_57_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _0911_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4014_ dacArea_dac_cnt_1\[0\] net63 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_84_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5965_ _1701_ _1702_ _1700_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4233__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4916_ dspArea_regB\[4\] _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5896_ _1198_ _3333_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5981__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4847_ _0696_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_14_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7566_ _0086_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5733__A2 _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4778_ _0272_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ _3490_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3729_ _3282_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7497_ _0017_ net217 dacArea_dac_cnt_5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _2281_ _2284_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5497__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6379_ _2209_ _2214_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_88_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5249__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6921__A1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__I dspArea_regB\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3840__I dspArea_regA\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ _1575_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6091__C _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _0554_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_37_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5681_ _1524_ _1453_ _1456_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7420_ _3225_ _3233_ _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4632_ _0440_ _0442_ _0439_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_8_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5715__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ dspArea_regP\[38\] _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4563_ dspArea_regP\[4\] _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6302_ _2027_ _2030_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7282_ _3055_ _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4494_ _0338_ _0357_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ _1962_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5007__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1901_ _1903_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _0954_ _0962_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _1934_ _1854_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6979__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _0892_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_2_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5651__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4206__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ _2721_ _2734_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_41_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ dspArea_regP\[20\] _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_80_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__A3 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5954__A2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5879_ _0989_ _1720_ _1721_ _1087_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6203__I0 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4509__A3 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7549_ _0069_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3925__I _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7506__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7395__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__I _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5945__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3835__I _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6211__I _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A2 _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4133__A1 _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _0349_ _3416_ _2662_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_39_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6851_ _2585_ _2682_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5802_ _1556_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3994_ dacArea_dac_cnt_0\[4\] net45 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6782_ _2550_ _2613_ _2615_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__5936__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _0514_ _3404_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7529__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _1276_ _1507_ _1508_ _1177_ _1285_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7403_ _3093_ _3220_ _3221_ _3224_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4615_ _0467_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3745__I dspArea_regA\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5595_ _1438_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__A1 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7334_ _3158_ _3118_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4546_ _0384_ _0385_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7265_ _3047_ _2454_ _3091_ _2855_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7310__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6216_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7196_ _3008_ _3023_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_48_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _1983_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _1879_ _1913_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0805_ _0878_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_45_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5927__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3938__A1 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7129__A1 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__S _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__I0 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6206__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ dspArea_regB\[2\] _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5380_ _0308_ _3346_ _1136_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ net101 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4106__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7050_ _2858_ _2879_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_87_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4262_ dacArea_dac_cnt_7\[3\] net55 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xfanout209 net223 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6001_ _1681_ _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5854__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__I _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4193_ dacArea_dac_cnt_5\[5\] net40 _3669_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_45_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5606__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6903_ _2721_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_82_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6834_ _2665_ _2666_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _0323_ _3443_ _2389_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3977_ _3489_ _3496_ _3497_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6582__A2 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7375__C _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _1539_ _1541_ _1558_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6696_ _2527_ _2530_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5647_ _1359_ _1378_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_40_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5578_ _1421_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input65_I user_clock2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _3119_ _3141_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4529_ _0386_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7248_ _3063_ _3074_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7179_ dspArea_regP\[34\] _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A3 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__A2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4820__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6573__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6325__A2 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5105__I dspArea_regA\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 la_data_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_37_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6261__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3900_ dspArea_regP\[18\] _3429_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4880_ _0662_ _0716_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _3374_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5775__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3762_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6550_ _2382_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5501_ _1345_ _1346_ _1145_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6481_ _2313_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5432_ _1274_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _1208_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _2920_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _0209_ _0204_ _0210_ _0206_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _0623_ _1039_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XDSP48_229 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5827__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4245_ dacArea_dac_cnt_7\[0\] net52 _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7033_ _2860_ _2861_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_19_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4176_ _3655_ _3654_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6252__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _2508_ _2567_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6555__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6748_ _2494_ _2495_ _2492_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_17_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6679_ _1233_ _2110_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3933__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5818__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__A3 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6491__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6243__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6546__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3843__I _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5809__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ dacArea_dac_cnt_1\[3\] net3 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5285__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6234__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1623_ _1714_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_64_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _0780_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7651_ net197 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4863_ _0713_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__A1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ _2343_ _2346_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_60_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3814_ _3359_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7582_ _0102_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__C _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4794_ _0603_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3756__C1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _2366_ _2367_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_21_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3745_ dspArea_regA\[1\] _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _2299_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5415_ _1157_ _1160_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3753__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _2068_ _2231_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xoutput132 net132 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput143 net143 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput154 net154 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4720__A1 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput165 net165 wb_DAT_MISO[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5346_ _0353_ _0501_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput176 net176 wb_DAT_MISO[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 net187 wb_DAT_MISO[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5277_ _1107_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6473__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ _2840_ _2843_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_4228_ dacArea_dac_cnt_6\[4\] net48 _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_75_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input28_I la_data_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ _3642_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5028__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5267__A2 dspArea_regA\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6767__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6415__S _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4778__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__B _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7192__A2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 la_data_in[1] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xinput23 la_data_in[2] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput34 la_data_in[3] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7562__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput45 la_data_in[4] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout215_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput56 la_data_in[5] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput67 wb_ADR[10] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 wb_ADR[20] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput89 wb_ADR[30] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5200_ _1042_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4702__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _2016_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _0898_ _0876_ _0979_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _0832_ _0844_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_69_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4013_ dacArea_dac_cnt_1\[0\] net63 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _1701_ _1702_ _1700_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_52_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _0755_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3748__I _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5895_ _1735_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4846_ dspArea_regP\[9\] _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5194__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _0085_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _3345_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _2045_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4941__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3728_ net91 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7496_ _0016_ net213 dacArea_dac_cnt_5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6447_ _2282_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5497__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6378_ _2115_ _2117_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6794__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _1082_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_87_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6446__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6997__A2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7585__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5185__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4932__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4489__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6685__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4160__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6437__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ dspArea_regA\[2\] _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3974__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5680_ _1357_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7165__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4631_ _0459_ _0484_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6912__A2 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ dspArea_regP\[37\] _3145_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4923__A1 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _0364_ _0420_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__A4 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _2048_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_7_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _3056_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4493_ _0356_ net104 _0344_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ _1967_ _1972_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4151__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ dspArea_regP\[21\] _1902_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _0851_ _0853_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7458__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _1840_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6979__A2 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5100__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5045_ _0893_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _2825_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__A2 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _0263_ _3447_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5878_ dspArea_regP\[19\] _1085_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I wb_ADR[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6203__I1 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5167__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4829_ _0297_ _3322_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__A2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4914__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ _0068_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7479_ _0153_ net207 dacArea_dac_cnt_3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6667__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3941__I _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__S _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__B _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A2 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__I dspArea_regA\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7600__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3851__I _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3892__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6850_ _2587_ _2588_ _2602_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1628_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _2460_ _2540_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3993_ _3499_ _3510_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_62_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5732_ _0623_ _3396_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _1174_ _1274_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7402_ _3194_ _3222_ _3223_ _3213_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__6897__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4614_ _0470_ _3314_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _1109_ dspArea_regA\[6\] _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7333_ _3104_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4372__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4545_ dspArea_regP\[2\] _0383_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7264_ _0988_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4476_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7310__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _1946_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7233__I _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _3012_ _3022_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5872__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _1984_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _1916_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6821__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _0805_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I la_data_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _0320_ _3465_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3936__I _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7408__I _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4115__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4666__A3 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6812__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__I dspArea_regB\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6415__I1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4426__I0 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A3 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4007__I _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6879__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _0221_ _0216_ _0222_ _0218_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_5_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5303__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _0164_ _0168_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _1671_ _1682_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_45_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _3667_ _3668_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input2_I la_data_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5606__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _2726_ _2731_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_36_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__I dspArea_regB\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__C _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _1755_ _3456_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A2 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _2595_ _2596_ _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3976_ _3494_ _3495_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5715_ _1539_ _1541_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__4593__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _2415_ _2528_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5646_ _1374_ _1377_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5542__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5577_ _1415_ _1417_ _1420_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7316_ _3122_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4528_ _0375_ _0376_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I la_data_in[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7247_ _3065_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4459_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7178_ _3001_ _3005_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _1968_ _3391_ _1756_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4281__A1 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4033__A1 _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__C2 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5881__I _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4497__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7519__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6261__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6013__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3830_ dspArea_regA\[11\] _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5772__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3761_ _3312_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5500_ _3390_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6480_ _2315_ _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _1276_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5524__A1 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5791__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _0330_ _0920_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7277__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7101_ _2928_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _3340_ _0201_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5293_ _1129_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7032_ _2813_ _2815_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5827__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4244_ dacArea_dac_cnt_7\[0\] net52 _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4175_ dacArea_dac_cnt_5\[1\] net36 _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input112_I wb_DAT_MOSI[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__A1 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _2508_ _2567_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4015__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _2579_ _2580_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3959_ dspArea_regP\[27\] _3486_ net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6678_ _2509_ _2512_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_52_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5629_ _0276_ _3403_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5515__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output164_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7440__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__A2 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A1 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5754__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5809__A2 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout195_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7491__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__S _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7431__A1 _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__A2 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5980_ _1616_ _1613_ _1715_ _1610_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _0693_ _0781_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7650_ net198 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4862_ _0603_ _0647_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6601_ _2359_ _2433_ _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3813_ _3358_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7581_ _0101_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4548__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _0643_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3756__B1 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6532_ _1636_ _3386_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3756__C2 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3744_ _3298_ net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6463_ _0607_ _3425_ _2199_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5414_ _1242_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _2131_ _2134_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput133 net133 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput144 net144 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0349_ _0501_ _1112_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput155 net155 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4720__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput166 net166 wb_DAT_MISO[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput177 net177 wb_DAT_MISO[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput188 net188 wb_DAT_MISO[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _1113_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7015_ _2844_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4227_ _3692_ _3696_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6473__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _3640_ _3637_ _3641_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_56_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7422__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _3491_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5984__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__A1 dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__A1 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput13 la_data_in[20] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput24 la_data_in[30] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput35 la_data_in[40] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput46 la_data_in[50] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput57 la_data_in[60] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3854__I dspArea_regA\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput68 wb_ADR[11] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__I _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput79 wb_ADR[21] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout208_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4702__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5130_ _0898_ _0876_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6455__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _0837_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_38_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ _3522_ _3526_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5963_ _1767_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _0759_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5894_ _1732_ _1733_ _1734_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_80_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _0697_ dspArea_regA\[9\] _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5718__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7564_ _0084_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4776_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _2348_ _2351_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3727_ net88 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7495_ _0015_ net216 dacArea_dac_cnt_5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6446_ _1323_ _1676_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6143__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ dspArea_regP\[23\] _2116_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5328_ _0994_ _0981_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input40_I la_data_in[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6446__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5259_ _1105_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A3 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6315__I _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5185__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6134__A1 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6685__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4630_ _0431_ _0485_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6373__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5176__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6912__A3 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4561_ dspArea_regP\[3\] _0419_ _0396_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4923__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _2052_ _2135_ _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7280_ _3070_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6125__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _0355_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6231_ _1967_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6676__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _1999_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A2 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5113_ dspArea_regP\[11\] _0852_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _1843_ _1853_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _0806_ _0803_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5100__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3759__I _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _0361_ _3410_ _2755_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_53_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ _1149_ _3439_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5877_ _1715_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _0607_ _3305_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6364__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input88_I wb_ADR[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7547_ _0067_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4759_ _0611_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4914__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6116__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7478_ _0152_ net207 dacArea_dac_cnt_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6667__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _1845_ _3378_ _2176_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_68_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6419__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7552__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4850__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4905__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5800_ _1631_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6780_ _2536_ _2539_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3992_ dacArea_dac_cnt_0\[4\] net45 _3509_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_50_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _1564_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6346__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _1282_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7401_ _3200_ _3214_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6897__A2 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5593_ _1437_ _3328_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7332_ _3099_ _3103_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4544_ _0399_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7263_ _3086_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6649__A2 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _1405_ _3348_ _1947_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7194_ _3014_ _3021_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _1352_ _3422_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7575__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6076_ _1782_ _1799_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5085__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4873__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6821__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _0806_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4832__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6978_ _1970_ _3457_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_81_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _0285_ _3425_ _1578_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6337__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5209__I dspArea_regA\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6812__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4823__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A1 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__I1 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A3 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6879__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7598__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ dacArea_dac_cnt_7\[3\] net55 _0167_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_5_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4191_ dacArea_dac_cnt_5\[4\] net39 _3664_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_45_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5789__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4814__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6901_ _2597_ _2732_ _2667_ _2664_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6832_ _0736_ _3448_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3975_ _3494_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6763_ _0314_ _3449_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4042__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6319__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _1543_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6694_ _2422_ _2423_ _2421_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5790__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ _1471_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5576_ _1415_ _1417_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_4527_ dspArea_regP\[1\] _0374_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7315_ _3139_ _3133_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3772__I _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7246_ _3071_ _3072_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4458_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7177_ _3003_ _3004_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4389_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _0320_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6059_ _1896_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_74_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3947__I dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5781__A2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3792__A1 dspArea_regP\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__B2 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5297__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6993__I _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4272__A2 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3857__I _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4024__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ dspArea_regA\[3\] _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _1174_ _1178_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5524__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _0339_ dspArea_regA\[3\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7100_ _2250_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4312_ net120 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5292_ _1138_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7031_ _2813_ _2815_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_87_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4243_ _3491_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4174_ _3559_ _3653_ _3654_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_45_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4263__A2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input105_I wb_DAT_MOSI[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _2638_ _2647_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_23_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__A1 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _2513_ _2526_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3958_ dspArea_regP\[26\] _3486_ net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5763__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3889_ _3426_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6677_ _2510_ _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6712__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5515__A2 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _1244_ _3395_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input70_I wb_ADR[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5559_ _1402_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7229_ _2874_ _2999_ _0328_ _3482_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5754__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4301__I _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5690__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6234__A3 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6672__B _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4930_ _0700_ _0702_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7195__A1 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _0643_ _0646_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6600_ _2434_ _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3812_ dspArea_regA\[9\] _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7580_ _0100_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4792_ _0560_ _0644_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5745__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3756__A1 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3756__B2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3743_ dspArea_regP\[32\] _3281_ _3289_ _3294_ _3297_ dspArea_regP\[0\] _3298_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6531_ _1527_ _3386_ _2284_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_14_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _0828_ _3441_ _2100_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _1256_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6393_ _2131_ _2134_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput134 net134 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5344_ _1190_ _3316_ _1015_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
Xoutput145 net145 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput156 net156 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput167 net167 wb_DAT_MISO[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput178 net178 wb_DAT_MISO[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput189 net189 wb_DAT_MISO[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5275_ _1119_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ dacArea_dac_cnt_6\[4\] net48 _3695_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_7014_ _2744_ _2745_ _2758_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_56_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4157_ dacArea_dac_cnt_4\[5\] net31 _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7422__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _3522_ _3586_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4236__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5984__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6933__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _1533_ _3393_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7509__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7110__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 la_data_in[21] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput25 la_data_in[31] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput36 la_data_in[41] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput47 la_data_in[51] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput58 la_data_in[61] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput69 wb_ADR[12] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3910__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7101__A1 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3870__I _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _0843_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4011_ net199 net62 _3525_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5415__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _1800_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_18_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__A1 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _0761_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7168__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5893_ _1732_ _1733_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ _0263_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5718__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7563_ _0083_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4775_ _0625_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6514_ _2349_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3726_ _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7494_ _0014_ net212 dacArea_dac_cnt_5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6445_ _1437_ _1058_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6143__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6376_ _2211_ _2213_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6577__B _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5327_ _0982_ _1083_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5258_ _1036_ _1049_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA_input33_I la_data_in[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ dacArea_dac_cnt_6\[1\] net44 _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_5_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ dspArea_regA\[10\] _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5957__A2 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7481__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6685__A3 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__B _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5948__A2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__A1 dspArea_regP\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3865__I _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout220_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4560_ _0398_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6125__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6230_ _1972_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5884__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__I _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6161_ dspArea_regP\[22\] _2000_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0957_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6092_ _3558_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5636__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5043_ _0877_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _2824_ _2754_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6061__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1783_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5876_ _1716_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _0676_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3775__I _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__A1 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7546_ _0066_ clknet_3_3__leaf_wb_clk_i dspArea_regB\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4758_ _0291_ _3315_ _0567_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3709_ net124 _zz_1_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7477_ _0151_ net210 dacArea_dac_cnt_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4689_ _0498_ _0541_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4390__A4 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6428_ _1414_ _3392_ _2077_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _0604_ _1992_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A1 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3810__C2 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__A2 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5866__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5618__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5094__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__I _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ _3507_ _3505_ _3508_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _1572_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_15_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5661_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6346__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__A1 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _3167_ _3219_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4612_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5592_ dspArea_regB\[12\] _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7331_ _3147_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4543_ dspArea_regP\[3\] _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7262_ _3087_ _3044_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4474_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _2049_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7193_ _3019_ _3020_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _0839_ _3414_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _1914_ _1915_ _1798_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6282__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5085__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5026_ _0873_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _2804_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6585__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _1768_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6337__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5859_ _1575_ _1593_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4348__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ _0049_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A2 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A3 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4304__I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6879__A3 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5000__A2 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ dacArea_dac_cnt_5\[4\] net39 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__A1 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4814__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _0323_ _3459_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _0928_ _3440_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A2 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _1450_ _2493_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ dacArea_dac_cnt_0\[1\] net12 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_17_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5713_ _1548_ _1553_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_6693_ _2422_ _2423_ _2421_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6319__A2 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ _1485_ _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5575_ _1419_ _3316_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7314_ _3138_ _3131_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7542__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4526_ _0384_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_2_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7245_ _0360_ _3452_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4457_ dspArea_regB\[10\] _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7176_ _2945_ _2950_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4388_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4884__I _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ _1963_ _1966_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _1897_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4805__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _0777_ _0779_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__A1 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6246__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4034__I _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7565__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4980__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _1011_ _0555_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4311_ _0207_ _0204_ _0208_ _0206_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ _1130_ _1131_ _1137_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6485__A1 dspArea_regP\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5288__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ _2808_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4242_ _3645_ _3708_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _3651_ _3652_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5460__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _2643_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6745_ _2578_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3957_ dspArea_regP\[25\] _3486_ net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6676_ _2417_ _2420_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3888_ _3425_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5627_ _0768_ _1059_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3783__I _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _1300_ _1313_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input63_I la_data_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _0267_ _3294_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_5489_ _1332_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6476__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5279__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7228_ _3051_ _3054_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_28_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _2986_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6228__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7588__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5203__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6467__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__I _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _0669_ _0709_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_72_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3811_ _3357_ net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _0577_ _0580_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_18_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6530_ _1632_ _3400_ _2175_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__3756__A2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3742_ _3296_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4699__I dspArea_regB\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _2296_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5412_ _1148_ _1257_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6392_ _2166_ _2226_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _0342_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput135 net135 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput146 net146 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput157 net157 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput168 net168 wb_DAT_MISO[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput179 net179 wb_DAT_MISO[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _1120_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_7013_ _2750_ _2757_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4225_ _3693_ _3690_ _3694_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ dacArea_dac_cnt_4\[5\] net31 _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ net197 net16 _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_55_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5433__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3778__I dspArea_regA\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A2 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4989_ _0839_ _0478_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ _2560_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6659_ _0924_ _2493_ _2288_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6697__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4402__I _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7110__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__I _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6924__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput15 la_data_in[22] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput26 la_data_in[32] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput37 la_data_in[42] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput48 la_data_in[52] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput59 la_data_in[62] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4312__I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7603__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ _3523_ _3519_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_78_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _1683_ _1801_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _0762_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _0353_ _3339_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_80_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7168__A2 _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _0694_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7562_ _0082_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4926__A1 dspArea_regP\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _0626_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6513_ _2239_ _2251_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3725_ net91 _3275_ _3279_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7493_ _0013_ net212 dacArea_dac_cnt_5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4222__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6679__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6444_ _1435_ _3384_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6375_ dspArea_regP\[24\] _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5326_ _1088_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _1042_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6851__A1 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ _3558_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _0950_ _0952_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input26_I la_data_in[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _3623_ _3626_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__I _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4145__A2 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5645__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout192 net151 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__I _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3959__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout213_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4977__I _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3881__I _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _1367_ dspArea_regA\[22\] _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5111_ dspArea_regP\[12\] _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _1830_ _0424_ _1931_ _1087_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5042_ _0888_ _0889_ _0890_ _0891_ _0795_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7389__A2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4447__I0 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6993_ _2753_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6061__A2 dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _1784_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_81_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ _1717_ _1617_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_61_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _0678_ _3324_ _0628_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4375__A2 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7545_ _0065_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _0547_ _0521_ _0517_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _0150_ net205 dacArea_dac_cnt_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4688_ _0497_ _0543_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _2263_ _2186_ _2189_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3791__I _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A2 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ _1886_ _3424_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_1_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _1148_ _1154_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6289_ _2005_ _2009_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A4 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A1 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7585__D _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3966__I _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__B2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7001__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5563__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7068__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5618__A2 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6517__I _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ dacArea_dac_cnt_0\[3\] net34 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _1392_ _1395_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ dspArea_regB\[2\] _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5554__A1 dspArea_regP\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4357__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5591_ _1435_ _3322_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7330_ _3152_ _3154_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4542_ _0266_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7261_ _3033_ _3036_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4473_ dspArea_regB\[12\] _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6212_ _2050_ _1950_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _1519_ _3444_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_48_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _1886_ _3407_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _1787_ _1794_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _0874_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_6_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7471__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A1 dacArea_dac_cnt_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6976_ _2805_ _2806_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ _0608_ _1229_ _1678_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_22_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3786__I dspArea_regA\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _1589_ _1592_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input93_I wb_ADR[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4348__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _0601_ _0602_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5789_ _0915_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7528_ _0048_ clknet_3_7__leaf_wb_clk_i dspArea_regA\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7459_ _0133_ net201 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5506__I _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4410__I _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A2 dspArea_regA\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4284__A1 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A3 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7289__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4320__I _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6264__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6830_ _2659_ _2662_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_63_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _1968_ _3441_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3973_ _3492_ _3493_ _3494_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _1554_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6692_ _2513_ _2526_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5643_ _1365_ _1486_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5574_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7313_ _3127_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4525_ _0274_ _3302_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7244_ _3069_ _3070_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _0311_ _0324_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7175_ _2941_ _3002_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6126_ _1964_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A3 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _1144_ _3438_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_74_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5008_ _0777_ _0779_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A2 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _2743_ _2759_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6191__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5236__I _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7443__A1 dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6067__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4980__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6182__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5146__I _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4310_ _3333_ _0201_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ _1130_ _1131_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ net193 net51 _3707_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6485__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4172_ _3651_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7434__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6237__A2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6813_ _2572_ _2644_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3956_ _3297_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6744_ _2510_ _2511_ _2509_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_52_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ dspArea_regP\[26\] _2416_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3887_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5626_ _1460_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5557_ _1303_ _1312_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4508_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _1333_ _0521_ _1215_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input56_I la_data_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__I dspArea_regB\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _3052_ _3053_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4439_ _0309_ net121 _0293_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7158_ _2888_ _2900_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_58_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _1947_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6228__A2 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7089_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4135__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6164__A1 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5911__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6467__A2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7181__I _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7416__A1 dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5978__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7532__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3810_ dspArea_regP\[40\] _3351_ _3342_ _3356_ _3349_ dspArea_regP\[8\] _3357_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_61_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _0577_ _0580_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3741_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3884__I dspArea_regA\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6460_ _2276_ _2278_ _2295_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6155__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5411_ _1154_ _1156_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6391_ _2092_ _2227_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5902__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5342_ _1187_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_12_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput136 net136 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput147 net147 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput158 net158 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput169 net169 wb_DAT_MISO[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5273_ _1019_ _0670_ _1024_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_7012_ _2842_ _2790_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ dacArea_dac_cnt_6\[3\] net47 _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5130__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4155_ _3622_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _3583_ _3581_ _3584_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5969__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__C _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input110_I wb_DAT_MOSI[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _0300_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_23_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6727_ _2557_ _2558_ _2559_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3939_ _3470_ _3471_ net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _3432_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _1434_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6589_ _2415_ _2421_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_3_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output162_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7555__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3969__I _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 la_data_in[23] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 la_data_in[33] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_6_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput38 la_data_in[43] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput49 la_data_in[53] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6688__A2 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5360__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout193_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3879__I _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5960_ _1696_ _1699_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4623__A1 dspArea_regP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _0297_ _0478_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5891_ _1416_ _3339_ _1654_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_61_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _3352_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ _0081_ clknet_3_1__leaf_wb_clk_i dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4926__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ _0277_ _3335_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3724_ net88 _3278_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6512_ _2235_ _2238_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7492_ _0012_ net211 dacArea_dac_cnt_5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6679__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6443_ _2193_ _2279_ _2202_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6374_ _0476_ dspArea_regA\[24\] _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ _1089_ _1170_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__7578__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _1048_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _3587_ _3679_ _3680_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_29_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _1034_ _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_5_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ dacArea_dac_cnt_4\[2\] net28 _3625_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3789__I _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I la_data_in[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ dacArea_dac_cnt_2\[3\] net11 _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4614__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6119__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout193 net150 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4081__A2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4323__I _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__B _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout206_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5333__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6530__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__I0 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5154__I _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _0477_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _1831_ _1929_ _1930_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6694__B _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _0806_ _0877_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__A2 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _2819_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_81_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4447__I1 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _0469_ _3431_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _1606_ _1609_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4825_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7544_ _0064_ clknet_3_1__leaf_wb_clk_i dspArea_regB\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5572__A2 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _0606_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5773__B _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7475_ _0149_ net204 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4687_ dspArea_regP\[6\] _0542_ _0396_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _2104_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6357_ _1348_ _3442_ _2112_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _1057_ _1061_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _2106_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0989_ _1084_ _1086_ _1087_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_76_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5260__A1 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__A2 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__A1 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7068__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5079__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4053__I _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _0465_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5590_ dspArea_regB\[13\] _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5554__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _3314_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7260_ _3037_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4472_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6211_ _1938_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7191_ _3017_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7059__A2 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6142_ _1348_ _3425_ _1899_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6073_ _1787_ _1794_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _0740_ _0793_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5490__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__B _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6034__A3 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6975_ _1110_ _2108_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4045__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ _0829_ _3399_ _1569_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _1683_ _1696_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4808_ _0660_ _0652_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5545__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ _1630_ _1557_ _1560_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input86_I wb_ADR[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _0047_ clknet_3_6__leaf_wb_clk_i dspArea_regA\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4739_ dspArea_regP\[7\] _0593_ _0396_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7458_ _0132_ net201 dacArea_dac_cnt_0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6409_ _1396_ _1504_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7389_ _3184_ _3187_ _3211_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6618__I dspArea_regP\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5522__I dspArea_regA\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7222__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5233__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5784__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__A1 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__A3 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4275__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5472__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4027__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3887__I _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6760_ _2590_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_50_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3972_ dacArea_dac_cnt_0\[0\] net1 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6972__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5711_ _1333_ _3346_ _1447_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6691_ _2517_ _2525_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5642_ _1371_ _1373_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6724__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ dspArea_regB\[14\] _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7312_ dspArea_regP\[37\] _1085_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4524_ dspArea_regP\[2\] _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7243_ _3066_ _3067_ _3068_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4455_ _0323_ net123 _0316_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7174_ _2944_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4386_ _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6125_ _1445_ _1676_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_58_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6056_ _0514_ _3431_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _0772_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__I _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6958_ _2743_ _2759_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_41_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _1749_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6889_ _2643_ _2646_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5252__I _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7443__A2 dspArea_regP\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A2 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4009__A2 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6182__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4331__I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7461__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _3705_ _3703_ _3706_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6485__A3 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A1 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4171_ dacArea_dac_cnt_5\[1\] net36 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5162__I dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__A1 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6812_ _2523_ _2640_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6743_ _2508_ _2567_ _2576_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_50_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3955_ _3484_ _3485_ net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _2507_ _2508_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3886_ _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5625_ _1468_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5556_ _1296_ _1391_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ _3271_ _3286_ _0366_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_5487_ _0747_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7226_ _0334_ _3480_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5684__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I la_data_in[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _2891_ _2899_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_8_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ _0240_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _1424_ _3348_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7088_ _2912_ _2916_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6039_ _1225_ _3408_ _1677_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4416__I _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5739__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7484__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7113__A1 _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _3282_ net91 _3275_ _3278_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_60_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6155__A2 dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4166__A1 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _1154_ _1156_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6390_ _2128_ _2129_ _2127_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5902__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5341_ _1103_ _1125_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7104__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput137 net137 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput148 net148 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput159 net159 wb_ACK vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5272_ _0737_ _3330_ _0921_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5666__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7011_ _2841_ _2742_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4223_ dacArea_dac_cnt_6\[3\] net47 _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4154_ _3623_ _3638_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4085_ dacArea_dac_cnt_2\[6\] net15 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input103_I wb_DAT_MOSI[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6394__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _0306_ _3323_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6726_ _2557_ _2558_ _2559_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3938_ dspArea_regP\[22\] _3463_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6657_ _2488_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3869_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5608_ _1441_ _1448_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_6588_ _2422_ _2423_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_11_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5539_ _1262_ _1263_ _1261_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7215__C _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7209_ _3033_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 la_data_in[24] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput28 la_data_in[34] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput39 la_data_in[44] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4623__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4910_ _0301_ _3323_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ _1190_ _3355_ _1546_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ dspArea_regB\[1\] _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__I dspArea_regA\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _0080_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4772_ _0515_ _3329_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _2256_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3723_ _3276_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7491_ _0011_ net213 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6442_ _2194_ _2195_ _2200_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6373_ _1150_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5324_ _1002_ _1078_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5639__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5255_ _1101_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6300__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__A3 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ dacArea_dac_cnt_6\[0\] net43 _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _0942_ _0945_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _3624_ _3621_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6064__A1 dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _3515_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6367__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A1 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _2543_ _2451_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6119__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7522__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4550__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4302__A1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout194 net148 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6055__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6358__A2 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7307__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6530__A2 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__I1 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7650__I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5097__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _0806_ _0877_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5170__I _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6046__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _2820_ _2821_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5942_ _0564_ _3423_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_46_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5873_ _1606_ _1609_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _0622_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ _0063_ clknet_3_5__leaf_wb_clk_i dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ _0608_ _3290_ _0557_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_30_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7545__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4780__A1 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5773__C _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7474_ _0148_ net206 dacArea_dac_cnt_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4686_ _0498_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6425_ _2095_ _2105_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__A1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ _1345_ _3458_ _1995_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ dspArea_regP\[13\] _1060_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6287_ _2122_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6285__A1 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5238_ _0240_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input31_I la_data_in[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5169_ dspArea_regB\[10\] _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5260__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4424__I _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4771__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__A2 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__A1 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6276__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7568__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _0274_ _3307_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4762__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4471_ _3487_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6210_ _1941_ _1949_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7190_ _1847_ _3452_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _1345_ _3442_ _1785_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1895_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _0789_ _0792_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6019__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6974_ _0996_ _3439_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ _1765_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6990__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _1581_ _1697_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4807_ _0545_ _0653_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_22_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5787_ _1469_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7526_ _0046_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4738_ _0544_ _0590_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA_input79_I wb_ADR[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7457_ _0131_ net200 dacArea_dac_cnt_0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4669_ _0273_ _3331_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4505__A1 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _2242_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7388_ _3173_ _3188_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6339_ _2173_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6258__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4419__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__A3 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6430__A1 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6249__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3971_ dacArea_dac_cnt_0\[0\] net1 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6972__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5710_ _0322_ _3360_ _1329_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6690_ _2521_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_52_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _1371_ _1373_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6724__A2 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _1416_ _3316_ _1325_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _0451_ _3135_ _3136_ _2855_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _0266_ _3307_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_7_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6488__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _3066_ _3067_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _2999_ _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6719__I _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ dspArea_regB\[0\] _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6124_ _1443_ _1058_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _0623_ _1582_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _0850_ _0854_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_73_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6957_ _2777_ _2780_ _2787_ _2786_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ _1110_ _0949_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4974__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6888_ _2718_ _2672_ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _1680_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4726__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7509_ _0029_ net218 dacArea_dac_cnt_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6479__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6651__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4593__B _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__B _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4612__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4193__A2 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6890__A1 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _3587_ _3650_ _3651_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3898__I _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6811_ _2569_ _2573_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6742_ _2571_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_56_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4956__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ dspArea_regP\[24\] _3463_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6673_ _2453_ _2504_ _2506_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_56_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3885_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4708__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5624_ _1461_ _1462_ _1467_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7370__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5555_ _1387_ _1390_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ net125 _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _0322_ _0631_ _1117_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _1413_ _3474_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4437_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5684__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7156_ _2980_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4368_ _3452_ _0247_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _1945_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7087_ _2912_ _2916_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ net117 _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _1877_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7229__B _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6787__C _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__A2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__I0 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6094__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3989__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__A2 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__A2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7653__I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ _1107_ _1124_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput127 net127 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput138 net138 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput149 net149 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5271_ _1114_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5173__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7010_ _2737_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4222_ _3622_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4153_ dacArea_dac_cnt_4\[5\] net31 _3637_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__5418__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ dacArea_dac_cnt_2\[6\] net15 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6091__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4986_ _0770_ _0833_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _3469_ _3453_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6725_ _1418_ _3400_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6656_ _2489_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3868_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _1449_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4157__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _2318_ _2325_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3799_ _3346_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5538_ _1262_ _1263_ _1261_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_3_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input61_I la_data_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _1219_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7208_ _3034_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6854__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _2859_ _2878_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_output148_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5593__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4162__I _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 la_data_in[25] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput29 la_data_in[35] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4148__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5345__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5896__A2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7098__A1 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4840_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4771_ _0624_ _3323_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6510_ _2259_ _2343_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3722_ net93 net95 net94 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7490_ _0010_ net213 dacArea_dac_cnt_4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6441_ _2177_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _3472_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5323_ _1074_ _1077_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5254_ _1017_ _1029_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4205_ dacArea_dac_cnt_6\[0\] net43 _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5185_ _1033_ _3346_ _0841_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_9_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ dacArea_dac_cnt_4\[1\] net27 _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7474__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6064__A2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4067_ _3543_ _3569_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_44_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5811__A2 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A2 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5575__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _0667_ _0816_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5078__I _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _2437_ _2440_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _1197_ _3387_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5878__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6827__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout195 net147 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6055__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A1 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6372__I _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7307__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__I _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__I _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6046__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _2717_ _2736_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5941_ _0562_ _3415_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7378__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5872_ _1623_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4823_ _0675_ _3338_ _0566_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_21_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7542_ _0062_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4754_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ _0147_ net206 dacArea_dac_cnt_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4685_ _0538_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4780__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6424_ _2161_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6355_ _2191_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4532__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6809__A1 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _1151_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6286_ _1998_ _2123_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6285__A2 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5237_ dspArea_regP\[13\] _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _1014_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_57_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input24_I la_data_in[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ dacArea_dac_cnt_3\[5\] net22 _3610_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__A1 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ dspArea_regA\[9\] _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4523__A2 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6276__A2 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A2 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4762__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout211_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _0311_ _0336_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7661__I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6140_ _1978_ _1979_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6071_ _1907_ _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5022_ _0808_ _0869_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6019__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A3 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _0347_ _2493_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_81_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _1743_ _1745_ _1764_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7512__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5855_ _1586_ _1588_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _0597_ _0656_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5786_ _1460_ _1470_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7525_ _0045_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4737_ _0591_ _0538_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5950__A1 dspArea_regP\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7456_ _0130_ net200 dacArea_dac_cnt_0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4668_ _0475_ _0480_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4505__A2 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _2048_ _2139_ _2241_ _2037_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5702__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ _3203_ _3209_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4599_ _0454_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _2174_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_143_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6258__A2 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6269_ _3447_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6915__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A2 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__I _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7446__A1 dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7535__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4680__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ _3491_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5640_ _1477_ _1482_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_31_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6724__A3 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5571_ _1305_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5932__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _0373_ _0377_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7310_ dspArea_regP\[36\] _0380_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_8_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6488__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _0354_ _3460_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4453_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7172_ _0328_ _3481_ _2869_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4384_ _0163_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7437__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6123_ _0927_ _3384_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_8_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _1882_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5999__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _0774_ _0776_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A2 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4671__A1 dspArea_regP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input126_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__I _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _2785_ _2770_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _0995_ _3352_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4974__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _2668_ _2671_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ _1672_ _1673_ _1679_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input91_I wb_ADR[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4726__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _1392_ _1395_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7508_ _0028_ net219 dacArea_dac_cnt_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6479__A2 dspArea_regA\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ dspArea_regP\[44\] _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7428__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__C _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__A2 dspArea_regA\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5914__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4717__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5390__A2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7419__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__A2 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3861__C1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _2639_ _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _2506_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3953_ _3483_ _3289_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_51_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6672_ _2504_ _2506_ _2453_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3884_ dspArea_regA\[17\] _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5905__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _1461_ _1462_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5554_ dspArea_regP\[17\] _0799_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_8_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4505_ net98 net159 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5485_ _1327_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7224_ _0350_ _3469_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4436_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6330__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ _2982_ _2983_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4367_ _0215_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5684__A3 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _1942_ _1943_ _1944_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7086_ _2913_ _2915_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _0197_ _0190_ _0198_ _0194_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_58_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6633__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6037_ _1857_ _1859_ _1876_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4644__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__C1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6397__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _2767_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_41_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6149__A1 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6321__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6872__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__I _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4635__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4486__I1 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5454__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput128 net128 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput139 net139 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _1115_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ _3666_ _3691_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4152_ _3635_ _3636_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4083_ _3570_ _3582_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6379__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7040__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4985_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6724_ _1527_ _3400_ _2486_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_51_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3936_ _3468_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6655_ _1116_ dspArea_regA\[19\] _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _3406_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5606_ _1450_ _3337_ _1330_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6551__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6586_ _2321_ _2324_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3798_ _3345_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5537_ _1340_ _1379_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5468_ _1300_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input54_I la_data_in[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7207_ _2985_ _2988_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4419_ _0268_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6854__A2 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5399_ _1144_ dspArea_regA\[13\] _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7103__I0 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7138_ _2862_ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7069_ _2897_ _2898_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5593__A2 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 la_data_in[26] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5345__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6542__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4084__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4353__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4770_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_61_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ net92 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6440_ _2182_ _2185_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6371_ _2205_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5184__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5322_ _1099_ _1166_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6836__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5253_ _1025_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4847__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _3645_ _3678_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5184_ _0302_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _3622_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ dacArea_dac_cnt_2\[3\] net11 _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_83_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A2 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A2 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4968_ _0814_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ _2457_ _2541_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3919_ _3452_ _3453_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4899_ _0739_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _2471_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6524__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _2207_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6827__A2 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4438__I _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout196 net146 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5978__B _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4066__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6515__A1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5318__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5940_ _1770_ _1781_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5871_ _1626_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _0284_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6754__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5557__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7541_ _0061_ clknet_3_2__leaf_wb_clk_i dspArea_regB\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4753_ _0551_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7472_ _0146_ net205 dacArea_dac_cnt_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5309__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ _0453_ _0492_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6423_ _1407_ _3363_ _2162_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6354_ _1342_ _1884_ _2101_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5305_ dspArea_regP\[14\] _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6285_ _2002_ _2004_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5236_ _0379_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5167_ _0997_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7591__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _3609_ _3607_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ _0937_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_17_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4048__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I la_data_in[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4049_ _3522_ _3555_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__I _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6200__A3 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7464__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout204_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5711__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _1908_ _1909_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4278__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I la_data_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5021_ _0752_ _0870_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6019__A3 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _2708_ _2709_ _2712_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6975__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5923_ _1743_ _1745_ _1764_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_80_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5854_ _1586_ _1588_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4805_ _0451_ _0657_ _0658_ _0261_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_10_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5785_ _1531_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7524_ _0044_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4736_ _0453_ _0492_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3961__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7455_ _0129_ net202 dacArea_dac_cnt_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4667_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6406_ _2141_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7386_ _3205_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5702__A2 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _0292_ _3292_ _0428_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6337_ _0331_ _1058_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_27_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6268_ _0624_ _3440_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5219_ _0954_ _1066_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _1816_ _1817_ _1928_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A1 dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__I _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5941__A2 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7143__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6249__A3 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ _1414_ _3332_ _1209_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5932__A2 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _0364_ _0381_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7672__I net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7240_ _2893_ _3460_ _2998_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4452_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _2995_ _2998_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4383_ _0259_ _0191_ _0260_ _0261_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5192__I _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _1958_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _1892_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5004_ dspArea_regP\[10\] _0775_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A3 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input119_I wb_DAT_MOSI[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _2785_ _2770_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_54_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5620__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5906_ _1012_ _0631_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6886_ _2663_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ _1672_ _1673_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_22_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5768_ _1296_ _1391_ _1503_ _1400_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4726__A3 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input84_I wb_ADR[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7507_ _0027_ net217 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4719_ _0571_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7125__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5699_ _1460_ _1542_ _1469_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7438_ _0369_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7369_ _3189_ _3192_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7428__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4111__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4662__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__A1 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A1 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7116__A1 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3861__B1 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3861__C2 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _2569_ _2572_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3952_ _3482_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6671_ _2404_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7355__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3883_ _3419_ _3421_ net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5622_ _1463_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_31_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5553_ _0882_ _1398_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4504_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5484_ _1328_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5669__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ dspArea_regP\[34\] _3006_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4435_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__A1 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7154_ _2884_ _2901_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_8_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4366_ net111 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _1942_ _1943_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_86_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _2914_ _2846_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4297_ _3308_ _0191_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _1857_ _1859_ _1876_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_55_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4644__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3852__B1 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__C2 dspArea_regP\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6397__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6938_ _2636_ _2768_ _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7346__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6869_ _2700_ _2701_ _2615_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6149__A2 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7525__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6321__A2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__I _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4635__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 dspArea_regB\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4946__I0 dspArea_regP\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4571__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput129 net129 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ dacArea_dac_cnt_6\[3\] net47 _3690_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ dacArea_dac_cnt_4\[4\] net30 _3633_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ dacArea_dac_cnt_2\[6\] net15 _3581_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5823__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6379__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _0465_ _0470_ _0834_ _0631_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6723_ _0334_ _3416_ _2467_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3935_ _3467_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7328__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7548__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6654_ _0735_ dspArea_regA\[18\] _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3866_ _3405_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6000__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ _0926_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6585_ _2417_ _2420_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_3797_ _3344_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4562__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _1380_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5467_ _1303_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7206_ _2980_ _2984_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4418_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5398_ _1244_ _0958_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input47_I la_data_in[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7137_ _2860_ _2861_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4349_ _0234_ _0227_ _0236_ _0229_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7103__I1 _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7068_ _1519_ _3427_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_28_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5814__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _1771_ _1772_ _1778_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_27_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5290__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7319__A1 dspArea_regP\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6790__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A2 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7098__A3 _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3803__I _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__A1 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _3271_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_13_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6370_ _2206_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_6_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5321_ _1032_ _1167_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_6_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5252_ _1028_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ net194 net42 _3677_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5183_ _1006_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _3488_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ dacArea_dac_cnt_2\[2\] net10 _3567_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5272__A2 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input101_I wb_DAT_MOSI[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6221__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ _0816_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3918_ _3310_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6706_ _2460_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4783__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4898_ _0746_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6637_ _2468_ _2469_ _2470_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3849_ _3390_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6524__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ _2403_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3743__C1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5519_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _2204_ _2221_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_65_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout197 net145 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__C _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4454__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6451__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5870_ _1709_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _0672_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7540_ _0060_ clknet_3_6__leaf_wb_clk_i dspArea_regA\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4752_ _0504_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4765__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7471_ _0145_ net203 dacArea_dac_cnt_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4683_ _0488_ _0491_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5309__A3 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _2257_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _1225_ _3433_ _1985_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5304_ _0476_ _3395_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6284_ _2002_ _2004_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5235_ _0991_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_88_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6690__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5166_ _0332_ _3304_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_64_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ dacArea_dac_cnt_3\[5\] net22 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _0941_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5245__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6442__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ net198 net7 _3554_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_25_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _1736_ _1839_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ net195 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5833__I dspArea_regA\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3731__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4449__I dspArea_regB\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6681__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6672__A1 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5475__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _0786_ _0787_ _0785_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _2799_ _2800_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_80_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6975__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4986__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5922_ _1747_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ _1689_ _1693_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ dspArea_regP\[8\] _0495_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4822__I _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5784_ _1406_ _3317_ _1532_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7523_ _0043_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4735_ _0545_ _0586_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_7454_ _0128_ net202 dacArea_dac_cnt_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3961__A2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4666_ dspArea_regP\[5\] _0265_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _2048_ _2139_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_7385_ _3206_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4597_ _0286_ _3307_ _0407_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_66_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6336_ _0995_ _3383_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4910__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6267_ _2095_ _2105_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5218_ _0962_ _0964_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ _0824_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__A2 _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7143__A2 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6654__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5393__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ dspArea_regP\[1\] _0378_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7581__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7170_ _2996_ _2997_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4382_ _0240_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__I _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6121_ _1959_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6645__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _1883_ _1885_ _1891_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__B _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5003_ _0851_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4120__A2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__A2 _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _2767_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5905_ _1671_ _1746_ _1681_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _2714_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5836_ _1674_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_14_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5384__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _1396_ _1504_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7506_ _0026_ net219 dacArea_dac_cnt_6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4718_ dspArea_regP\[7\] _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_5698_ _1461_ _1462_ _1467_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input77_I wb_ADR[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7437_ _3225_ _3244_ _3253_ _3254_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4649_ _0303_ _3291_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _3190_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _1413_ _3386_ _1960_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7299_ _3063_ _3074_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7454__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5611__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__A2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__I _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__A1 dspArea_regP\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3861__B2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3951_ _3481_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _0561_ _3478_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3882_ dspArea_regP\[16\] _3420_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1464_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5366__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5552_ dspArea_regP\[16\] _1397_ _0726_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4503_ _3274_ _3284_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5483_ _1022_ _1045_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5669__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7222_ _3029_ _3032_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4434_ dspArea_regB\[7\] _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7153_ _2981_ _2883_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4365_ _0246_ _0238_ _0248_ _0241_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _1419_ _3355_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _2840_ _2843_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7477__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ net116 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _1861_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5841__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A1 dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__B2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6937_ _2693_ _2696_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_41_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4282__I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _2630_ _2631_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7346__A2 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5819_ _1450_ _0834_ _1552_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6799_ _2609_ _2612_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6203__S _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output183_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4457__I dspArea_regB\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4096__A1 _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A2 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7034__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__I1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4571__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5520__A1 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ dacArea_dac_cnt_4\[4\] net30 _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7273__A1 dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__I _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ dacArea_dac_cnt_2\[5\] net14 _3580_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__A1 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _0695_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _2555_ _2497_ _2500_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3934_ _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7328__A2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _1018_ _3423_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3865_ _3404_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5604_ _0924_ _0834_ _1214_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4011__A1 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6584_ _2403_ _2418_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3796_ _3343_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5535_ _1242_ _1260_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6839__A1 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5466_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7205_ _3029_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4417_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5511__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ dspArea_regB\[3\] _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7136_ _2963_ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4348_ _3410_ _0235_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7264__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ _2895_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _0181_ _0179_ _0182_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4078__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5814__A2 dspArea_regA\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6018_ _1752_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4250__A1 _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A2 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5571__I _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6616__B _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5741__A1 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5320_ _1071_ _1072_ _1070_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_6_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6297__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _1092_ _1098_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4202_ _3675_ _3673_ _3676_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1010_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_9_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4133_ _3559_ _3620_ _3621_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_60_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4064_ _3564_ _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_7_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7515__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6221__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4232__A1 _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _0313_ _3312_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6705_ _2536_ _2539_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3917_ _3451_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5980__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0748_ _3290_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _2468_ _2469_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_22_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6524__A3 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5732__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _0464_ _3472_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3779_ _3328_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3743__B1 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3743__C2 dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5518_ _1360_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6498_ _2217_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_79_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5449_ _1186_ _1294_ _1293_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__3904__I _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output146_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _0333_ _3466_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_87_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout198 net144 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7267__B _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4774__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5971__A1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3814__I _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7538__CLK clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A2 dspArea_regA\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7400__A1 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _0309_ _0501_ _0618_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4751_ _0604_ _0555_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4380__I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7470_ _0144_ net205 dacArea_dac_cnt_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4682_ _0499_ _0534_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6421_ _2153_ _2165_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4517__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6352_ _2188_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _1150_ _3390_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6283_ _2114_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _0994_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_9_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7219__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _1013_ _0552_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4116_ _3596_ _3608_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _0942_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4555__I _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4047_ _3552_ _3550_ _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6442__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1407_ _3333_ _1737_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5953__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ dspArea_regP\[11\] _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5386__I dspArea_regB\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4290__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ net196 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ _0422_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5705__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7599_ _0119_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A2 _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4465__I _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__A2 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5296__I dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3809__I _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7449__A1 dspArea_regP\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4683__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _2731_ _2733_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _1752_ _1758_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_34_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ _1583_ _1585_ _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _0597_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_61_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5783_ _1624_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7522_ _0042_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4734_ _0499_ _0587_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7453_ _0127_ net202 dacArea_dac_cnt_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4665_ _3329_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6404_ _1821_ _1822_ _2039_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7384_ _3175_ _3183_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_31_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6360__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _0445_ _0444_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6335_ _1012_ _3376_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _2103_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4486__S _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6663__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _0962_ _0964_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6197_ _2034_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5148_ _0996_ _3299_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input22_I la_data_in[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4285__I _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _0928_ _0461_ _0818_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__A2 dspArea_regA\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4450_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6342__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4381_ _3483_ _0189_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6893__A2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ _1323_ _3374_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6645__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _1883_ _1885_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__C _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ dspArea_regP\[11\] _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_78_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7070__A2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ dspArea_regP\[31\] _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _1672_ _1673_ _1679_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6884_ _2638_ _2647_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5908__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5835_ _1675_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ _1606_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__4187__A3 _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6581__A1 dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5384__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7505_ _0025_ net219 dacArea_dac_cnt_6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4717_ _0477_ _3344_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5697_ _1441_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ dspArea_regP\[43\] _3365_ _3238_ _3245_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ _0298_ _3300_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6333__A1 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7367_ _3161_ _3165_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4579_ dspArea_regP\[3\] _0401_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6318_ _2155_ _2088_ _2091_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7298_ _3065_ _3073_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6249_ _2079_ _2084_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__3912__I dspArea_regA\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6572__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5574__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__A2 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__I _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3861__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _3411_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5620_ _0554_ _3383_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5366__A2 dspArea_regA\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5551_ _1292_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _0337_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5482_ _0319_ _0689_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7221_ _3024_ _3028_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4433_ _0288_ _0304_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4877__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7152_ _2880_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4364_ _3444_ _0247_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _1416_ _3355_ _1865_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _2840_ _2843_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4295_ _0195_ _0190_ _0196_ _0194_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _1866_ _1871_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__C1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input124_I wb_STB vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__I dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _2693_ _2696_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_70_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _2630_ _2631_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_23_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ _0924_ _3367_ _1446_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6798_ _2613_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5749_ _1589_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__3907__I _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7419_ _3229_ _3232_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6953__I dspArea_regP\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7571__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A2 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__I _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__I dspArea_regB\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__A2 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3817__I _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__I _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _3579_ _3577_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4087__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4982_ _0756_ _0771_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6721_ _2413_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3933_ _3465_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _2484_ _2486_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5339__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ _3403_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__I0 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _1442_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6583_ _0278_ _3478_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4011__A2 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3727__I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3795_ dspArea_regA\[7\] _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5534_ _1256_ _1259_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6839__A2 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5465_ _1197_ _3301_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7204_ _3030_ _3031_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4416_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5511__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _0768_ _3375_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7135_ _2897_ _2898_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4347_ _0200_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7594__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7264__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7066_ _0354_ _3435_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4278_ dacArea_dac_cnt_7\[6\] net59 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5275__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _1758_ _1762_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4293__I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6919_ _1632_ _3434_ _2592_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6527__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4561__I0 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4468__I _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6616__C _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6766__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6518__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7191__A1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _1096_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ dacArea_dac_cnt_5\[6\] net41 _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_64_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _1017_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4132_ _3618_ _3619_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5257__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4063_ dacArea_dac_cnt_2\[2\] net10 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6757__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A3 _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4965_ _0815_ dspArea_regA\[2\] _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6704_ _2375_ _2537_ _2538_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4841__I dspArea_regB\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _3450_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5980__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _0352_ _3392_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3847_ dspArea_regA\[13\] _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _2400_ _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3778_ dspArea_regA\[5\] _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5732__A2 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3743__A1 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _1361_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3743__B2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ _2219_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__I _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _1189_ _1201_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input52_I la_data_in[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4288__I _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5379_ _1225_ _3361_ _1046_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _0915_ _3458_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xfanout199 net143 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7049_ _2859_ _2863_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_41_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7267__C _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3830__I dspArea_regA\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5411__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ _0300_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5962__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3973__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7164__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _0459_ _0535_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_18_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _2156_ _2164_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5714__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6351_ _2168_ _2170_ _2187_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5302_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6282_ _2118_ _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3740__A4 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5478__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5233_ _1079_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__7413__S _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4115_ dacArea_dac_cnt_3\[5\] net22 _3607_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__4836__I _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _0943_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4046_ dacArea_dac_cnt_1\[6\] net6 _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6442__A3 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4205__A2 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _1836_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4948_ _0370_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7667_ net197 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _0713_ _0715_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_14_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6618_ dspArea_regP\[27\] _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7598_ _0118_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6549_ _2383_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3915__I _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__I dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5944__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__A1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7146__A1 _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3825__I _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7505__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4683__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5880__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _1760_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ dspArea_regP\[18\] _1584_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__I _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4199__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _0652_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5782_ _1522_ _1536_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_15_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7521_ _0041_ clknet_3_2__leaf_wb_clk_i dspArea_regA\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4733_ _0534_ _0537_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7452_ _0126_ net202 dacArea_dac_cnt_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4664_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6403_ _2031_ _2140_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_31_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7383_ dspArea_regP\[38\] _3174_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4595_ _0446_ _0444_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3735__I dspArea_regA\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6334_ _2095_ _2171_ _2104_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6265_ _2096_ _2097_ _2102_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5216_ _1056_ _1062_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6196_ _1813_ _1815_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_57_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5871__A1 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4566__I _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5147_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I la_data_in[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ dacArea_dac_cnt_1\[3\] net3 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5397__I dspArea_regB\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__A2 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7528__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4901__A3 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6103__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4476__I _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3928__A1 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7119__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6342__A2 _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout202_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4380_ net115 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6866__I _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1887_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I la_data_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4386__I _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _0477_ _3375_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6952_ _1932_ _2783_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_19_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _1655_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6883_ dspArea_regP\[29\] _2637_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _0295_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5908__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3919__A1 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5765_ _1404_ _1607_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5384__A3 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4592__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7504_ _0024_ net219 dacArea_dac_cnt_6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4716_ _0570_ _3338_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5696_ _1448_ _1452_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7435_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4647_ _0500_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6333__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__A1 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _3156_ _3160_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4578_ _0432_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_11_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ _1989_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7297_ _3119_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _2085_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_76_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4296__I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _1879_ _2017_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_58_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6021__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6572__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__I dspArea_regB\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _3417_ _3418_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_56_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4574__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _1392_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_12_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _0338_ _0363_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5481_ _0927_ _0769_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7220_ dspArea_regP\[35\] _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4326__A1 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ _0303_ net120 _0293_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _2961_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4363_ _0188_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1190_ _3370_ _1750_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7082_ _2907_ _2911_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _3302_ _0191_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A1 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _1872_ _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__B1 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__C2 dspArea_regP\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4844__I _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7220__I dspArea_regP\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6251__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input117_I wb_DAT_MOSI[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _2763_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_42_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _2616_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6003__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5817_ _1656_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5675__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6797_ _2550_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _1477_ _1590_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input82_I wb_ADR[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _1344_ _1358_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_11_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__A1 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ _3237_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _3152_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__3923__I _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4754__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5808__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6481__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__I _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _0830_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6784__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ dspArea_regA\[22\] _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6720_ _2402_ _2414_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _2467_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3863_ dspArea_regA\[15\] _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6536__A2 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5602_ _1444_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4398__I1 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ _0622_ _2314_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3794_ _3288_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5533_ _1359_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _1308_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7203_ _2965_ _2978_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4415_ dspArea_regB\[4\] _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5395_ _1228_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7134_ _2962_ _2896_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4346_ net105 _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _2892_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4277_ dacArea_dac_cnt_7\[6\] net59 _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_41_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _1758_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5275__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__A2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _2747_ _2748_ _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6849_ _2587_ _2588_ _2602_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3918__I _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4710__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A2 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4484__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6766__A2 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4241__A3 _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3828__I _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4529__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ dacArea_dac_cnt_5\[6\] net41 _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5180_ _1025_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _3618_ _3619_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ _3543_ _3565_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4394__I dspArea_regB\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4964_ _0318_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6703_ _2429_ _2432_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3915_ _3449_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3738__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ dspArea_regB\[10\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3846_ _3388_ net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6634_ _1305_ _3392_ _2385_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3777_ _3327_ net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6565_ _0760_ _3433_ _2307_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_69_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7561__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3743__A2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ _0276_ dspArea_regA\[14\] _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6496_ _2113_ _2121_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5447_ _1189_ _1201_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5378_ _0302_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input45_I la_data_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7117_ _1634_ _3451_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4329_ _3371_ _0212_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6445__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7048_ _2868_ _2873_ _2877_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6684__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5239__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4998__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6739__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5411__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7584__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _0484_ _0487_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_41_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _2168_ _2170_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4922__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ dspArea_regB\[1\] _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4389__I _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ _1999_ _2001_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5478__A2 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6675__A1 dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _1080_ _0993_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4150__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5163_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_9_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4114_ _3605_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5094_ _0296_ _0689_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6978__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ dacArea_dac_cnt_1\[6\] net6 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4989__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ _1728_ _1740_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _0497_ _0798_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_33_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4461__I0 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ net198 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _0719_ _0717_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_71_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6617_ _2355_ _0424_ _2452_ _2354_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5166__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ _3288_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5683__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _0117_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _0330_ dspArea_regA\[15\] _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_3_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4299__I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _0469_ dspArea_regA\[23\] _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output151_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7457__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6969__A2 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7218__I0 dspArea_regP\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4904__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3841__I _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6409__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5850_ _1690_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _0545_ _0653_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__A1 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1525_ _1535_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7520_ _0040_ clknet_3_3__leaf_wb_clk_i dspArea_regA\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _0534_ _0537_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5148__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7451_ _0125_ clknet_3_0__leaf_wb_clk_i _zz_1_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4663_ _0513_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6402_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6896__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7382_ dspArea_regP\[39\] _3204_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4594_ _0426_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6333_ _2096_ _2097_ _2102_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6648__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _2096_ _2097_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _0957_ _0961_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4123__A2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3751__I dspArea_regA\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _1725_ _1833_ _1834_ _1927_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _0339_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3882__A1 dspArea_regP\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5077_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6820__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4028_ _3516_ _3538_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__I _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5979_ _1819_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5926__A3 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7128__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7649_ net199 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3926__I _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6887__A1 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__A3 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4492__I _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7119__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0570_ _3368_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ dspArea_regP\[30\] _2782_ _2628_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _1660_ _1663_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6882_ dspArea_regP\[30\] _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_34_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ dspArea_regA\[14\] _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _1499_ _1502_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7503_ _0023_ net216 dacArea_dac_cnt_6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4715_ _0272_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5695_ _1448_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7434_ dspArea_regP\[43\] dspArea_regP\[42\] _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4646_ _0292_ _0501_ _0472_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6333__A3 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _3173_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4577_ dspArea_regP\[4\] _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_2_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _1980_ _1990_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7296_ _3120_ _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _1970_ _3385_ _1966_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5844__A2 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6178_ _1916_ _1917_ _1913_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7046__A1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _0901_ _0905_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_45_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__A1 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6021__A2 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5835__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4271__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4023__A1 _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4500_ _0362_ net105 _0344_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5480_ _1321_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_144_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4431_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5523__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ _2965_ _2978_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4362_ net109 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4397__I _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1940_ _1875_ _1878_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6079__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7081_ _2910_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4293_ net110 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _1333_ _3368_ _1757_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__A1 dspArea_regP\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3837__B2 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A1 dspArea_regP\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7518__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6251__A2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6934_ _2764_ _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _2633_ _2697_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6003__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1657_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _1932_ _2629_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_10_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5747_ _1482_ _1484_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5762__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input75_I wb_ADR[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7417_ dspArea_regP\[41\] _3236_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5514__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0436_ _0438_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7348_ _3154_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7267__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7279_ _3071_ _3072_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__I _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4005__A1 _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5505__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5106__I _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7430__A1 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4980_ _0608_ _0400_ _0764_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_17_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3931_ _3462_ _3464_ net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_16_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _1323_ _1368_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3862_ _3402_ net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5601_ _1445_ dspArea_regA\[9\] _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4547__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ dspArea_regP\[26\] _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3793_ _3341_ net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5532_ _1374_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ _1304_ _1306_ _1307_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7202_ _2970_ _2977_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4414_ _0163_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5394_ _1239_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7133_ _2895_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4345_ _0232_ _0227_ _0233_ _0229_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4276_ _0164_ _0180_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7064_ _2893_ _3434_ _2807_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6472__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _1762_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7490__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _2658_ _2673_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4786__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6848_ _2561_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_50_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ _2609_ _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3934__I _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4710__A2 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7412__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6766__A3 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3844__I _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4130_ dacArea_dac_cnt_4\[1\] net27 _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4061_ dacArea_dac_cnt_2\[2\] net10 _3564_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__6454__A2 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _0327_ _0462_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6702_ _2429_ _2432_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3914_ _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ _0738_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_60_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _2283_ _2467_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3845_ dspArea_regP\[44\] _3382_ _3373_ _3387_ _3380_ dspArea_regP\[12\] _3388_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_34_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6564_ _0828_ _3450_ _2198_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6390__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3776_ dspArea_regP\[36\] _3320_ _3311_ _3326_ _3318_ dspArea_regP\[4\] _3327_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_9_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5515_ _1244_ _3389_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3754__I _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6495_ _2312_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6130__I _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6142__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5446_ _1287_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _1222_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7116_ _2941_ _2944_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4328_ net100 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input38_I la_data_in[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6445__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _2875_ _2876_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4259_ dacArea_dac_cnt_7\[2\] net54 _0166_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_47_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3929__I _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3982__A3 _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6133__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4998__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3839__I _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4922__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6124__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6280_ dspArea_regP\[22\] _2000_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5231_ _0974_ _0977_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5162_ dspArea_regB\[13\] _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ dacArea_dac_cnt_3\[4\] net21 _3603_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5093_ _0507_ _3336_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _3543_ _3551_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_37_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4989__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5650__A3 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5938__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _1731_ _1739_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_52_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4946_ dspArea_regP\[10\] _0797_ _0726_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4610__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__I1 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7665_ net199 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _0723_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6616_ _2450_ _2451_ _0367_ _0986_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_3828_ _3372_ net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5166__A2 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _0116_ clknet_3_3__leaf_wb_clk_i dspArea_regP\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6902__A3 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6547_ dspArea_regB\[12\] _1676_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3759_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6115__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _0464_ _2314_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_79_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6418__A2 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output144_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7091__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7218__I1 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6354__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__A2 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__CLK clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _0586_ _0589_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6593__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5396__A2 _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5780_ _1518_ _1621_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4731_ _0546_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _3489_ _3264_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4662_ _0516_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__6345__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _2235_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6896__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7381_ _0362_ _3483_ _3148_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0421_ _0424_ _0450_ _0261_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6332_ _2079_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_6_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6263_ _2098_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ dspArea_regP\[12\] _0960_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6194_ _1835_ _2032_ _2033_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5145_ _0901_ _0992_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__3882__A2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5076_ dspArea_regB\[10\] _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5084__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4027_ dacArea_dac_cnt_1\[3\] net3 _3537_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_38_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6820__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5978_ _1623_ _1714_ _1606_ _1609_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_12_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _0700_ _0702_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5694__I _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6336__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6887__A2 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7579_ _0099_ clknet_3_7__leaf_wb_clk_i dspArea_regP\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6639__A2 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__I _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A3 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__A2 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5075__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__A2 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6575__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6878__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5109__I _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5550__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4948__I _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5853__A3 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5066__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6950_ _2771_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _1660_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_19_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6881_ _2710_ _2712_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ dspArea_regB\[6\] _3389_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _1499_ _1502_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7502_ _0022_ net216 dacArea_dac_cnt_6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4714_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5694_ _1452_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7433_ _2856_ _3251_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4645_ _3300_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7364_ _3184_ _3187_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4576_ _0266_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6315_ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7295_ _3059_ _3075_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7597__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6246_ _1968_ _3398_ _1869_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_39_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6177_ _1916_ _1917_ _1913_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_58_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__A2 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0974_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA_input20_I la_data_in[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5057__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _0907_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__A1 dspArea_regP\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__A2 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6309__A1 _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4768__I dspArea_regB\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A2 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__A3 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7037__A2 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6548__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3847__I dspArea_regA\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4430_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6720__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4361_ _0244_ _0238_ _0245_ _0241_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_4_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _1780_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _2908_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4292_ _0185_ _0190_ _0192_ _0194_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _0322_ _3385_ _1658_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6933_ _2681_ _2691_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4262__A2 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6864_ _2636_ _2693_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_35_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A3 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ _1116_ dspArea_regA\[11\] _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_23_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6795_ dspArea_regP\[28\] _2627_ _2628_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3757__I _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5211__A1 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1482_ _1484_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5677_ _1422_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7416_ dspArea_regP\[41\] _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4628_ _0436_ _0438_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6711__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5514__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input68_I wb_ADR[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7347_ _3498_ _3137_ _3171_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_11_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _0413_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7267__A2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _3099_ _3103_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6229_ _2055_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_58_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4253__A2 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6043__I _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4498__I _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A1 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7430__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ dspArea_regP\[21\] _3463_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3861_ dspArea_regP\[46\] _3382_ _3373_ _3401_ _3380_ dspArea_regP\[14\] _3402_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_32_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5600_ dspArea_regB\[8\] _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6580_ dspArea_regP\[25\] _1150_ _3478_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_3792_ dspArea_regP\[38\] _3320_ _3311_ _3340_ _3318_ dspArea_regP\[6\] _3341_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ _1249_ _1375_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ _1304_ _1306_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7201_ _3024_ _3028_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4413_ _0262_ _0287_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_5393_ _1230_ _1231_ _1238_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7132_ _2957_ _2960_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _3401_ _0224_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7063_ _1634_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4275_ dacArea_dac_cnt_7\[6\] net59 _0179_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _1840_ _1854_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_39_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6472__A3 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5032__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input122_I wb_DAT_MOSI[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _2658_ _2673_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_35_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6847_ _0361_ _3393_ _2562_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_39_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6932__A1 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6778_ _2477_ _2610_ _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5735__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ _1565_ _1566_ _1571_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__A2 dspArea_regA\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__I _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A1 _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6923__A1 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__A2 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7508__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4537__I0 dspArea_regP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7100__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3860__I _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4060_ _3563_ _3562_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4962_ _0811_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _2477_ _2532_ _2535_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_3913_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7167__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ _0314_ _3304_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ dspArea_regB\[12\] _3403_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3844_ _3386_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6914__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _2397_ _2398_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3775_ _3325_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6390__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5514_ _0289_ _0959_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6494_ _2326_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5445_ _1288_ _1289_ _1290_ _1283_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6142__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6693__A3 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _1203_ _1204_ _1221_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3900__A1 dspArea_regP\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7115_ _2942_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_59_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4327_ _0219_ _0216_ _0220_ _0218_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3770__I dspArea_regA\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _0328_ _3459_ _2812_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4258_ _0161_ _0165_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4189_ _3622_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5405__A1 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7158__A1 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3719__A1 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6133__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4776__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A1 dspArea_regP\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__A1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout218_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7480__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6124__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _1002_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5161_ _1008_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_9_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4112_ dacArea_dac_cnt_3\[4\] net21 _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5092_ _0614_ _3330_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5635__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ dacArea_dac_cnt_1\[6\] net6 _3550_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_84_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _1725_ _1833_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_24_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6060__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _0729_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7664_ net192 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4876_ _0717_ _0720_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3827_ _3365_ _3351_ _3342_ _3371_ _3349_ dspArea_regP\[10\] _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_21_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6615_ _2447_ _2449_ _2441_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7595_ _0115_ clknet_3_0__leaf_wb_clk_i dspArea_regP\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3765__I _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7237__I _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6546_ _1011_ _1059_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ _3287_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7312__A1 dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ dspArea_regA\[22\] _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4126__A1 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _1088_ _1173_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input50_I la_data_in[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__A1 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ _1129_ _1205_ _1139_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _2706_ _2707_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_74_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7379__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5929__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6354__A2 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4500__S _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5617__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4730_ _0581_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _0468_ _3321_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__6345__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6400_ _2052_ _2236_ _2237_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_80_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7380_ _3178_ _3182_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4592_ _0426_ _0448_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _2084_ _2087_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_7_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _2099_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_66_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5213_ _1057_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6193_ _1838_ _2028_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4349__C _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5144_ _0905_ _0978_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_57_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6845__B _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5075_ _0924_ _3314_ _0745_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_56_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ dacArea_dac_cnt_1\[2\] net2 _3536_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6820__A3 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _1623_ _1714_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ _0772_ _0777_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input98_I wb_CYC vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6336__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _0710_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ _0098_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _2364_ _2294_ _2297_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7064__A3 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5838__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A1 dspArea_regP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__I _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5066__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5900_ _1663_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6880_ _2639_ _2642_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ dspArea_regB\[7\] _0959_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4577__A1 dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5762_ _1518_ _1602_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_7501_ _0021_ net216 dacArea_dac_cnt_6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4713_ _0563_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5693_ _1522_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4329__A1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7432_ dspArea_regP\[43\] _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_4644_ _0286_ _0400_ _0427_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6869__A3 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7363_ _3185_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4575_ _3321_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6314_ _2063_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_7294_ _3050_ _3058_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5829__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _2080_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _1977_ _2011_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_58_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5127_ _0827_ _0975_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7046__A3 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ _0335_ _0390_ _0823_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_73_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I la_data_in[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ dacArea_dac_cnt_0\[6\] net61 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7541__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A2 dspArea_regA\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3863__I dspArea_regA\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout200_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _3435_ _0235_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _0193_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _1867_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I la_data_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6932_ _2684_ _2690_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4643__B _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6863_ _2566_ _2694_ _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _0735_ dspArea_regA\[10\] _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_22_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6794_ _0395_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5211__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1581_ _1586_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_13_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7564__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ _1519_ _3308_ _1423_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7415_ dspArea_regP\[40\] _3231_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_11_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4627_ _0474_ _0481_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _0799_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4558_ _0415_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7277_ dspArea_regP\[36\] _3102_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4489_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6475__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6228_ _2058_ _2066_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _0271_ _3456_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5202__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3749__C1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6466__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A2 dspArea_regA\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7430__A3 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__I _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3860_ _3400_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3791_ _3339_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _1253_ _1255_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5461_ _0352_ _3306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7200_ _3026_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4412_ _0286_ net117 _0269_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4704__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _1230_ _1231_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_7131_ _2958_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4343_ net104 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _0343_ _3451_ _2724_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_4274_ dacArea_dac_cnt_7\[5\] net58 _0178_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_59_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _1843_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_41_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A1 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input115_I wb_DAT_MOSI[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _2655_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3768__I _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _2677_ _2603_ _2678_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_51_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _2532_ _2535_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3989_ dacArea_dac_cnt_0\[3\] net34 _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6932__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _1565_ _1566_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA_input80_I wb_ADR[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ _1401_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_11_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7329_ _3113_ _3153_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_output167_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5671__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6687__A1 dspArea_regB\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__I1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7100__A2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__A1 dspArea_regP\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout198_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _0755_ _0766_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _2399_ _2533_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_51_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3912_ dspArea_regA\[20\] _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4892_ _0742_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _2465_ _2395_ _2398_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5178__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3843_ _3385_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6914__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3774_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6562_ _2377_ _2379_ _2396_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4640__C _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5513_ _1344_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6493_ _2327_ _2328_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_12_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5444_ _0982_ _1083_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7602__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4153__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _1203_ _1204_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7114_ _2871_ _2872_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4326_ _3363_ _0212_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4257_ dacArea_dac_cnt_7\[2\] net54 _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7045_ _2729_ _2874_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5043__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4188_ _3639_ _3665_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3967__A2 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6829_ _2660_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3719__A2 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7330__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__A3 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__A1 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4455__I0 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7149__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__A2 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7321__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__A1 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3871__I _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _0935_ _0936_ _0947_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4111_ _3596_ _3604_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_69_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5091_ _0847_ _0938_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_42_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ dacArea_dac_cnt_1\[5\] net5 _3549_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6832__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5399__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ _1810_ _1811_ _1809_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6060__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4944_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7663_ net193 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _0497_ _0727_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_36_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6614_ _2441_ _2447_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
X_3826_ _3370_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7594_ _0114_ clknet_3_6__leaf_wb_clk_i dspArea_regP\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6363__A3 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6545_ _2301_ _2380_ _2310_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3757_ _3309_ net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6476_ _0677_ _3457_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7312__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1184_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3781__I _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5874__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5358_ _1130_ _1131_ _1137_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input43_I la_data_in[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ net119 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5289_ _1132_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_59_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7028_ dspArea_regP\[32\] _2857_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_28_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7091__A4 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A3 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4062__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3956__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7000__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6354__A3 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4117__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5865__A2 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5617__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6290__A2 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3866__I _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4660_ _0515_ _3312_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__A3 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _0444_ _0447_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6330_ _2084_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_143_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4108__A2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__I dspArea_regA\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__A1 dspArea_regP\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _1775_ _1992_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5212_ dspArea_regP\[13\] _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1838_ _2028_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_5143_ _0905_ _0978_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__A1 dspArea_regP\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _0320_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4025_ _3533_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6417__I dspArea_regP\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _1816_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4595__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5792__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _0696_ _0699_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4858_ _0621_ _0642_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3809_ _3355_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7577_ _0097_ clknet_3_5__leaf_wb_clk_i dspArea_regP\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4789_ _0621_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_14_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6528_ _2202_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _2276_ _2278_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_69_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__I dspArea_regB\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5847__A2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A3 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4283__A1 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__A1 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _0290_ _3397_ _1579_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5761_ _1603_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7500_ _0020_ net214 dacArea_dac_cnt_6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _0565_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ _1525_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7431_ _0154_ _3249_ _3250_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ _0454_ _0455_ _0457_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5526__A1 dspArea_regP\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _3147_ _3155_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4574_ _0273_ _0400_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1405_ _3356_ _2064_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_144_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7293_ _3104_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__5829__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _2081_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ _2013_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5126_ _0866_ _0867_ _0863_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__A2 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _0819_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4008_ dacArea_dac_cnt_0\[6\] net61 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5765__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _1696_ _1699_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__C2 dspArea_regP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A3 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7442__A1 dspArea_regP\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__I _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__C2 dspArea_regP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4290_ net126 _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7433__A1 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6931_ _2743_ _2759_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_48_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6862_ _2606_ _2607_ _2604_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_34_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _0325_ _0949_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_62_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5747__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6795__I0 dspArea_regP\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _2616_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_22_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ _1479_ _1481_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _0359_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4970__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7414_ _2856_ _3235_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4626_ _0432_ _0435_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7345_ _3140_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4557_ _0280_ _3293_ _0389_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7276_ _3100_ _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4488_ dspArea_regB\[14\] _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__I _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6227_ _2064_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_77_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6089_ _1817_ _1832_ _1928_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3749__B1 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__A1 dspArea_regP\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6466__A2 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__A1 dspArea_regP\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ _3338_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3874__I dspArea_regA\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _1305_ _3306_ _1210_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__6154__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5901__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _1232_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_7130_ _2858_ _2879_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4342_ _0230_ _0227_ _0231_ _0229_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_67_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ _2889_ _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4273_ _0177_ _0175_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1851_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
.ends

